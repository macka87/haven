-- desc_man_pkg.vhd: Descriptor manager package
-- Copyright (C) 2006 CESNET
-- Author(s): Lukas Solanka <solanka@liberouter.org>
--
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above copyright
--    notice, this list of conditions and the following disclaimer in
--    the documentation and/or other materials provided with the
--    distribution.
-- 3. Neither the name of the Company nor the names of its contributors
--    may be used to endorse or promote products derived from this
--    software without specific prior written permission.
--
-- This software is provided ``as is'', and any express or implied
-- warranties, including, but not limited to, the implied warranties of
-- merchantability and fitness for a particular purpose are disclaimed.
-- In no event shall the company or contributors be liable for any
-- direct, indirect, incidental, special, exemplary, or consequential
-- damages (including, but not limited to, procurement of substitute
-- goods or services; loss of use, data, or profits; or business
-- interruption) however caused and on any theory of liability, whether
-- in contract, strict liability, or tort (including negligence or
-- otherwise) arising in any way out of the use of this software, even
-- if advised of the possibility of such damage.
--
-- $Id$
--
-- TODO:
--
--
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
use IEEE.std_logic_arith.all;

-- ----------------------------------------------------------------------------
--                        DESC_MAN Package
-- ----------------------------------------------------------------------------
package desc_man_pkg is
   
   -- Initialization detect bit position
   -- Change only this constant if you need it
   constant DESC_MAN_INIT_BIT_POS : integer := 18;

   -- Initialization offset based on INIT_BIT_POS
   constant DESC_MAN_INIT_PHASE_OFFSET : std_logic_vector(31 downto 0) :=
      conv_std_logic_vector(2**DESC_MAN_INIT_BIT_POS, 32);
   

end desc_man_pkg;


-- ----------------------------------------------------------------------------
--                        DESC_MAN Package
-- ----------------------------------------------------------------------------
package body desc_man_pkg is
       
end desc_man_pkg;

