-------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /    Vendor: Xilinx
-- \   \   \/     Version : 1.6
--  \   \         Application : RocketIO GTX Wizard
--  /   /         Filename : ROCKETIO_WRAPPER.vhd
-- /___/   /\     Timestamp : 02/08/2005 09:12:43
-- \   \  /  \
--  \___\/\___\
--
--
-- Module ROCKETIO_WRAPPER (a GTX Wrapper)
-- Generated by Xilinx RocketIO GTX Wizard

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;


--***************************** Entity Declaration ****************************

entity ROCKETIO_WRAPPER is
generic
(
    -- Simulation attributes
    WRAPPER_SIM_MODE                : string    := "FAST"; -- Set to Fast Functional Simulation Model
    WRAPPER_SIM_GTXRESET_SPEEDUP    : integer   := 0; -- Set to 1 to speed up sim reset
    WRAPPER_SIM_PLL_PERDIV2         : bit_vector:= x"140"; -- Set to the VCO Unit Interval time
    --
    CH01_SWAP   : boolean := false;     -- TRUE to swap XAUI channels 1 and 2
    CH23_SWAP   : boolean := false      -- TRUE to swap XAUI channels 3 and 4
);
port
(

    --_________________________________________________________________________
    --_________________________________________________________________________
    --TILE0  (Location)

    ------------------------ Loopback and Powerdown Ports ----------------------
    TILE0_LOOPBACK0_IN                      : in   std_logic_vector(2 downto 0);
    TILE0_LOOPBACK1_IN                      : in   std_logic_vector(2 downto 0);
    TILE0_RXPOWERDOWN0_IN                   : in   std_logic_vector(1 downto 0);
    TILE0_RXPOWERDOWN1_IN                   : in   std_logic_vector(1 downto 0);
    TILE0_TXPOWERDOWN0_IN                   : in   std_logic_vector(1 downto 0);
    TILE0_TXPOWERDOWN1_IN                   : in   std_logic_vector(1 downto 0);
    ----------------------- Receive Ports - 8b10b Decoder ----------------------
    TILE0_RXCHARISCOMMA0_OUT                : out  std_logic_vector(1 downto 0);
    TILE0_RXCHARISCOMMA1_OUT                : out  std_logic_vector(1 downto 0);
    TILE0_RXCHARISK0_OUT                    : out  std_logic_vector(1 downto 0);
    TILE0_RXCHARISK1_OUT                    : out  std_logic_vector(1 downto 0);
    TILE0_RXDISPERR0_OUT                    : out  std_logic_vector(1 downto 0);
    TILE0_RXDISPERR1_OUT                    : out  std_logic_vector(1 downto 0);
    TILE0_RXNOTINTABLE0_OUT                 : out  std_logic_vector(1 downto 0);
    TILE0_RXNOTINTABLE1_OUT                 : out  std_logic_vector(1 downto 0);
    ------------------- Receive Ports - Channel Bonding Ports ------------------
    TILE0_RXCHANBONDSEQ0_OUT                : out  std_logic;
    TILE0_RXCHANBONDSEQ1_OUT                : out  std_logic;
    TILE0_RXENCHANSYNC0_IN                  : in   std_logic;
    TILE0_RXENCHANSYNC1_IN                  : in   std_logic;
    ------------------- Receive Ports - Clock Correction Ports -----------------
    TILE0_RXCLKCORCNT0_OUT                  : out  std_logic_vector(2 downto 0);
    TILE0_RXCLKCORCNT1_OUT                  : out  std_logic_vector(2 downto 0);
    --------------- Receive Ports - Comma Detection and Alignment --------------
    TILE0_RXBYTEISALIGNED0_OUT              : out  std_logic;
    TILE0_RXBYTEISALIGNED1_OUT              : out  std_logic;
    TILE0_RXBYTEREALIGN0_OUT                : out  std_logic;
    TILE0_RXBYTEREALIGN1_OUT                : out  std_logic;
    TILE0_RXCOMMADET0_OUT                   : out  std_logic;
    TILE0_RXCOMMADET1_OUT                   : out  std_logic;
    TILE0_RXENMCOMMAALIGN0_IN               : in   std_logic;
    TILE0_RXENMCOMMAALIGN1_IN               : in   std_logic;
    TILE0_RXENPCOMMAALIGN0_IN               : in   std_logic;
    TILE0_RXENPCOMMAALIGN1_IN               : in   std_logic;
    ------------------- Receive Ports - RX Data Path interface -----------------
    TILE0_RXDATA0_OUT                       : out  std_logic_vector(15 downto 0);
    TILE0_RXDATA1_OUT                       : out  std_logic_vector(15 downto 0);
    TILE0_RXRESET0_IN                       : in   std_logic;
    TILE0_RXRESET1_IN                       : in   std_logic;
    TILE0_RXUSRCLK0_IN                      : in   std_logic;
    TILE0_RXUSRCLK1_IN                      : in   std_logic;
    TILE0_RXUSRCLK20_IN                     : in   std_logic;
    TILE0_RXUSRCLK21_IN                     : in   std_logic;
    ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    TILE0_RXCDRRESET0_IN                    : in   std_logic;
    TILE0_RXCDRRESET1_IN                    : in   std_logic;
    TILE0_RXELECIDLE0_OUT                   : out  std_logic;
    TILE0_RXELECIDLE1_OUT                   : out  std_logic;
    TILE0_RXN0_IN                           : in   std_logic;
    TILE0_RXN1_IN                           : in   std_logic;
    TILE0_RXP0_IN                           : in   std_logic;
    TILE0_RXP1_IN                           : in   std_logic;
    -------- Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
    TILE0_RXBUFRESET0_IN                    : in   std_logic;
    TILE0_RXBUFRESET1_IN                    : in   std_logic;
    TILE0_RXBUFSTATUS0_OUT                  : out  std_logic_vector(2 downto 0);
    TILE0_RXBUFSTATUS1_OUT                  : out  std_logic_vector(2 downto 0);
    TILE0_RXCHANISALIGNED0_OUT              : out  std_logic;
    TILE0_RXCHANISALIGNED1_OUT              : out  std_logic;
    TILE0_RXCHANREALIGN0_OUT                : out  std_logic;
    TILE0_RXCHANREALIGN1_OUT                : out  std_logic;
    --------------- Receive Ports - RX Loss-of-sync State Machine --------------
    TILE0_RXLOSSOFSYNC0_OUT                 : out  std_logic_vector(1 downto 0);
    TILE0_RXLOSSOFSYNC1_OUT                 : out  std_logic_vector(1 downto 0);
    -------------- Receive Ports - polarity  -----------------------------------
    TILE0_RXPOLARITY0                       : in   std_logic;
    TILE0_RXPOLARITY1                       : in   std_logic;
    ------------- Shared Ports - Dynamic Reconfiguration Port (DRP) ------------
    TILE0_DADDR_IN                          : in   std_logic_vector(6 downto 0);
    TILE0_DCLK_IN                           : in   std_logic;
    TILE0_DEN_IN                            : in   std_logic;
    TILE0_DI_IN                             : in   std_logic_vector(15 downto 0);
    TILE0_DO_OUT                            : out  std_logic_vector(15 downto 0);
    TILE0_DRDY_OUT                          : out  std_logic;
    TILE0_DWE_IN                            : in   std_logic;
    --------------------- Shared Ports - Tile and PLL Ports --------------------
    TILE0_CLKIN_IN                          : in   std_logic;
    TILE0_GTXRESET_IN                       : in   std_logic;
    TILE0_PLLLKDET_OUT                      : out  std_logic;
    TILE0_REFCLKOUT_OUT                     : out  std_logic;
    TILE0_RESETDONE0_OUT                    : out  std_logic;
    TILE0_RESETDONE1_OUT                    : out  std_logic;
    ---------------- Transmit Ports - 8b10b Encoder Control Ports --------------
    TILE0_TXCHARISK0_IN                     : in   std_logic_vector(1 downto 0);
    TILE0_TXCHARISK1_IN                     : in   std_logic_vector(1 downto 0);
    ------------------ Transmit Ports - TX Data Path interface -----------------
    TILE0_TXDATA0_IN                        : in   std_logic_vector(15 downto 0);
    TILE0_TXDATA1_IN                        : in   std_logic_vector(15 downto 0);
    TILE0_TXRESET0_IN                       : in   std_logic;
    TILE0_TXRESET1_IN                       : in   std_logic;
    TILE0_TXUSRCLK0_IN                      : in   std_logic;
    TILE0_TXUSRCLK1_IN                      : in   std_logic;
    TILE0_TXUSRCLK20_IN                     : in   std_logic;
    TILE0_TXUSRCLK21_IN                     : in   std_logic;
    --------------- Transmit Ports - TX Driver and OOB signalling --------------
    TILE0_TXN0_OUT                          : out  std_logic;
    TILE0_TXN1_OUT                          : out  std_logic;
    TILE0_TXP0_OUT                          : out  std_logic;
    TILE0_TXP1_OUT                          : out  std_logic;
    -------- Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
    TILE0_TXENPMAPHASEALIGN0_IN             : in   std_logic;
    TILE0_TXENPMAPHASEALIGN1_IN             : in   std_logic;
    TILE0_TXPMASETPHASE0_IN                 : in   std_logic;
    TILE0_TXPMASETPHASE1_IN                 : in   std_logic;
    -------------- Transmit Ports - polarity  ----------------------------------
    TILE0_TXPOLARITY0                       : in   std_logic;
    TILE0_TXPOLARITY1                       : in   std_logic;
    ----------------- Transmit Ports - TX Ports for PCI Express ----------------
    TILE0_TXELECIDLE0_IN                    : in   std_logic;
    TILE0_TXELECIDLE1_IN                    : in   std_logic;



    --_________________________________________________________________________
    --_________________________________________________________________________
    --TILE1  (Location)

    ------------------------ Loopback and Powerdown Ports ----------------------
    TILE1_LOOPBACK0_IN                      : in   std_logic_vector(2 downto 0);
    TILE1_LOOPBACK1_IN                      : in   std_logic_vector(2 downto 0);
    TILE1_RXPOWERDOWN0_IN                   : in   std_logic_vector(1 downto 0);
    TILE1_RXPOWERDOWN1_IN                   : in   std_logic_vector(1 downto 0);
    TILE1_TXPOWERDOWN0_IN                   : in   std_logic_vector(1 downto 0);
    TILE1_TXPOWERDOWN1_IN                   : in   std_logic_vector(1 downto 0);
    ----------------------- Receive Ports - 8b10b Decoder ----------------------
    TILE1_RXCHARISCOMMA0_OUT                : out  std_logic_vector(1 downto 0);
    TILE1_RXCHARISCOMMA1_OUT                : out  std_logic_vector(1 downto 0);
    TILE1_RXCHARISK0_OUT                    : out  std_logic_vector(1 downto 0);
    TILE1_RXCHARISK1_OUT                    : out  std_logic_vector(1 downto 0);
    TILE1_RXDISPERR0_OUT                    : out  std_logic_vector(1 downto 0);
    TILE1_RXDISPERR1_OUT                    : out  std_logic_vector(1 downto 0);
    TILE1_RXNOTINTABLE0_OUT                 : out  std_logic_vector(1 downto 0);
    TILE1_RXNOTINTABLE1_OUT                 : out  std_logic_vector(1 downto 0);
    ------------------- Receive Ports - Channel Bonding Ports ------------------
    TILE1_RXCHANBONDSEQ0_OUT                : out  std_logic;
    TILE1_RXCHANBONDSEQ1_OUT                : out  std_logic;
    TILE1_RXENCHANSYNC0_IN                  : in   std_logic;
    TILE1_RXENCHANSYNC1_IN                  : in   std_logic;
    ------------------- Receive Ports - Clock Correction Ports -----------------
    TILE1_RXCLKCORCNT0_OUT                  : out  std_logic_vector(2 downto 0);
    TILE1_RXCLKCORCNT1_OUT                  : out  std_logic_vector(2 downto 0);
    --------------- Receive Ports - Comma Detection and Alignment --------------
    TILE1_RXBYTEISALIGNED0_OUT              : out  std_logic;
    TILE1_RXBYTEISALIGNED1_OUT              : out  std_logic;
    TILE1_RXBYTEREALIGN0_OUT                : out  std_logic;
    TILE1_RXBYTEREALIGN1_OUT                : out  std_logic;
    TILE1_RXCOMMADET0_OUT                   : out  std_logic;
    TILE1_RXCOMMADET1_OUT                   : out  std_logic;
    TILE1_RXENMCOMMAALIGN0_IN               : in   std_logic;
    TILE1_RXENMCOMMAALIGN1_IN               : in   std_logic;
    TILE1_RXENPCOMMAALIGN0_IN               : in   std_logic;
    TILE1_RXENPCOMMAALIGN1_IN               : in   std_logic;
    ------------------- Receive Ports - RX Data Path interface -----------------
    TILE1_RXDATA0_OUT                       : out  std_logic_vector(15 downto 0);
    TILE1_RXDATA1_OUT                       : out  std_logic_vector(15 downto 0);
    TILE1_RXRESET0_IN                       : in   std_logic;
    TILE1_RXRESET1_IN                       : in   std_logic;
    TILE1_RXUSRCLK0_IN                      : in   std_logic;
    TILE1_RXUSRCLK1_IN                      : in   std_logic;
    TILE1_RXUSRCLK20_IN                     : in   std_logic;
    TILE1_RXUSRCLK21_IN                     : in   std_logic;
    ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    TILE1_RXCDRRESET0_IN                    : in   std_logic;
    TILE1_RXCDRRESET1_IN                    : in   std_logic;
    TILE1_RXELECIDLE0_OUT                   : out  std_logic;
    TILE1_RXELECIDLE1_OUT                   : out  std_logic;
    TILE1_RXN0_IN                           : in   std_logic;
    TILE1_RXN1_IN                           : in   std_logic;
    TILE1_RXP0_IN                           : in   std_logic;
    TILE1_RXP1_IN                           : in   std_logic;
    -------- Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
    TILE1_RXBUFRESET0_IN                    : in   std_logic;
    TILE1_RXBUFRESET1_IN                    : in   std_logic;
    TILE1_RXBUFSTATUS0_OUT                  : out  std_logic_vector(2 downto 0);
    TILE1_RXBUFSTATUS1_OUT                  : out  std_logic_vector(2 downto 0);
    TILE1_RXCHANISALIGNED0_OUT              : out  std_logic;
    TILE1_RXCHANISALIGNED1_OUT              : out  std_logic;
    TILE1_RXCHANREALIGN0_OUT                : out  std_logic;
    TILE1_RXCHANREALIGN1_OUT                : out  std_logic;
    --------------- Receive Ports - RX Loss-of-sync State Machine --------------
    TILE1_RXLOSSOFSYNC0_OUT                 : out  std_logic_vector(1 downto 0);
    TILE1_RXLOSSOFSYNC1_OUT                 : out  std_logic_vector(1 downto 0);
    -------------- Receive Ports - polarity  -----------------------------------
    TILE1_RXPOLARITY0                       : in   std_logic;
    TILE1_RXPOLARITY1                       : in   std_logic;
    ------------- Shared Ports - Dynamic Reconfiguration Port (DRP) ------------
    TILE1_DADDR_IN                          : in   std_logic_vector(6 downto 0);
    TILE1_DCLK_IN                           : in   std_logic;
    TILE1_DEN_IN                            : in   std_logic;
    TILE1_DI_IN                             : in   std_logic_vector(15 downto 0);
    TILE1_DO_OUT                            : out  std_logic_vector(15 downto 0);
    TILE1_DRDY_OUT                          : out  std_logic;
    TILE1_DWE_IN                            : in   std_logic;
    --------------------- Shared Ports - Tile and PLL Ports --------------------
    TILE1_CLKIN_IN                          : in   std_logic;
    TILE1_GTXRESET_IN                       : in   std_logic;
    TILE1_PLLLKDET_OUT                      : out  std_logic;
    TILE1_REFCLKOUT_OUT                     : out  std_logic;
    TILE1_RESETDONE0_OUT                    : out  std_logic;
    TILE1_RESETDONE1_OUT                    : out  std_logic;
    ---------------- Transmit Ports - 8b10b Encoder Control Ports --------------
    TILE1_TXCHARISK0_IN                     : in   std_logic_vector(1 downto 0);
    TILE1_TXCHARISK1_IN                     : in   std_logic_vector(1 downto 0);
    ------------------ Transmit Ports - TX Data Path interface -----------------
    TILE1_TXDATA0_IN                        : in   std_logic_vector(15 downto 0);
    TILE1_TXDATA1_IN                        : in   std_logic_vector(15 downto 0);
    TILE1_TXRESET0_IN                       : in   std_logic;
    TILE1_TXRESET1_IN                       : in   std_logic;
    TILE1_TXUSRCLK0_IN                      : in   std_logic;
    TILE1_TXUSRCLK1_IN                      : in   std_logic;
    TILE1_TXUSRCLK20_IN                     : in   std_logic;
    TILE1_TXUSRCLK21_IN                     : in   std_logic;
    --------------- Transmit Ports - TX Driver and OOB signalling --------------
    TILE1_TXN0_OUT                          : out  std_logic;
    TILE1_TXN1_OUT                          : out  std_logic;
    TILE1_TXP0_OUT                          : out  std_logic;
    TILE1_TXP1_OUT                          : out  std_logic;
    -------- Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
    TILE1_TXENPMAPHASEALIGN0_IN             : in   std_logic;
    TILE1_TXENPMAPHASEALIGN1_IN             : in   std_logic;
    TILE1_TXPMASETPHASE0_IN                 : in   std_logic;
    TILE1_TXPMASETPHASE1_IN                 : in   std_logic;
    -------------- Transmit Ports - polarity  ----------------------------------
    TILE1_TXPOLARITY0                       : in   std_logic;
    TILE1_TXPOLARITY1                       : in   std_logic;        
    ----------------- Transmit Ports - TX Ports for PCI Express ----------------
    TILE1_TXELECIDLE0_IN                    : in   std_logic;
    TILE1_TXELECIDLE1_IN                    : in   std_logic
);

    attribute X_CORE_INFO : string;
    attribute X_CORE_INFO of ROCKETIO_WRAPPER  : entity is "gtxwizard_v1_6, Coregen v11.2";
end ROCKETIO_WRAPPER;

architecture RTL of ROCKETIO_WRAPPER is

--***************************** Signal Declarations *****************************

    -- Channel Bonding Signals
    signal  tile0_rxchbondo0_i   : std_logic_vector(3 downto 0);
    signal  tile0_rxchbondo1_i   : std_logic_vector(3 downto 0);

    -- CC_2B_1SKP Signals
    signal  tile0_rxdata0_i                 : std_logic_vector(15 downto 0);
    signal  tile0_rxcharisk0_i              : std_logic_vector(1 downto 0);
    signal  tile0_rxchariscomma0_i          : std_logic_vector(1 downto 0);
    signal  tile0_rxrundisp0_i              : std_logic_vector(1 downto 0);
    signal  tile0_rxnotintable0_i           : std_logic_vector(1 downto 0);
    signal  tile0_rxdisperr0_i              : std_logic_vector(1 downto 0);
    signal  tile0_rxbufstatus0_i            : std_logic_vector(2 downto 0);
    signal  tile0_rxclkcorcnt0_i            : std_logic_vector(2 downto 0);
    signal  tile0_rxchanbondseq0_i          : std_logic;
    signal  tile0_rxchanisaligned0_i        : std_logic;
    signal  tile0_rxchanrealign0_i          : std_logic;
    signal  tile0_rxlossofsync0_i           : std_logic_vector(1 downto 0);
    signal  tile0_rxvalid0_i                : std_logic;
    signal  tile0_rxrecclk0_i               : std_logic;
    signal  tile0_resetdone0_i              : std_logic;
    signal  tile0_rxreset0_i                : std_logic;
    signal  tile0_rxbufreset0_i             : std_logic;
    signal  tile0_rxdata1_i                 : std_logic_vector(15 downto 0);
    signal  tile0_rxcharisk1_i              : std_logic_vector(1 downto 0);
    signal  tile0_rxchariscomma1_i          : std_logic_vector(1 downto 0);
    signal  tile0_rxrundisp1_i              : std_logic_vector(1 downto 0);
    signal  tile0_rxnotintable1_i           : std_logic_vector(1 downto 0);
    signal  tile0_rxdisperr1_i              : std_logic_vector(1 downto 0);
    signal  tile0_rxbufstatus1_i            : std_logic_vector(2 downto 0);
    signal  tile0_rxclkcorcnt1_i            : std_logic_vector(2 downto 0);
    signal  tile0_rxchanbondseq1_i          : std_logic;
    signal  tile0_rxchanisaligned1_i        : std_logic;
    signal  tile0_rxchanrealign1_i          : std_logic;
    signal  tile0_rxlossofsync1_i           : std_logic_vector(1 downto 0);
    signal  tile0_rxvalid1_i                : std_logic;
    signal  tile0_rxrecclk1_i               : std_logic;
    signal  tile0_resetdone1_i              : std_logic;
    signal  tile0_rxreset1_i                : std_logic;
    signal  tile0_rxbufreset1_i             : std_logic;


    signal  tile1_rxchbondo0_i   : std_logic_vector(3 downto 0);
    signal  tile1_rxchbondo1_i   : std_logic_vector(3 downto 0);

    -- CC_2B_1SKP Signals
    signal  tile1_rxdata0_i                 : std_logic_vector(15 downto 0);
    signal  tile1_rxcharisk0_i              : std_logic_vector(1 downto 0);
    signal  tile1_rxchariscomma0_i          : std_logic_vector(1 downto 0);
    signal  tile1_rxrundisp0_i              : std_logic_vector(1 downto 0);
    signal  tile1_rxnotintable0_i           : std_logic_vector(1 downto 0);
    signal  tile1_rxdisperr0_i              : std_logic_vector(1 downto 0);
    signal  tile1_rxbufstatus0_i            : std_logic_vector(2 downto 0);
    signal  tile1_rxclkcorcnt0_i            : std_logic_vector(2 downto 0);
    signal  tile1_rxchanbondseq0_i          : std_logic;
    signal  tile1_rxchanisaligned0_i        : std_logic;
    signal  tile1_rxchanrealign0_i          : std_logic;
    signal  tile1_rxlossofsync0_i           : std_logic_vector(1 downto 0);
    signal  tile1_rxvalid0_i                : std_logic;
    signal  tile1_rxrecclk0_i               : std_logic;
    signal  tile1_resetdone0_i              : std_logic;
    signal  tile1_gtp0_cc_2b_1skp_reset_i   : std_logic;
    signal  tile1_rxrecclk0_bufg_i          : std_logic;
    signal  tile1_rxreset0_i                : std_logic;
    signal  tile1_rxbufreset0_i             : std_logic;
    signal  tile1_rxdata1_i                 : std_logic_vector(15 downto 0);
    signal  tile1_rxcharisk1_i              : std_logic_vector(1 downto 0);
    signal  tile1_rxchariscomma1_i          : std_logic_vector(1 downto 0);
    signal  tile1_rxrundisp1_i              : std_logic_vector(1 downto 0);
    signal  tile1_rxnotintable1_i           : std_logic_vector(1 downto 0);
    signal  tile1_rxdisperr1_i              : std_logic_vector(1 downto 0);
    signal  tile1_rxbufstatus1_i            : std_logic_vector(2 downto 0);
    signal  tile1_rxclkcorcnt1_i            : std_logic_vector(2 downto 0);
    signal  tile1_rxchanbondseq1_i          : std_logic;
    signal  tile1_rxchanisaligned1_i        : std_logic;
    signal  tile1_rxchanrealign1_i          : std_logic;
    signal  tile1_rxlossofsync1_i           : std_logic_vector(1 downto 0);
    signal  tile1_rxvalid1_i                : std_logic;
    signal  tile1_rxrecclk1_i               : std_logic;
    signal  tile1_resetdone1_i              : std_logic;
    signal  tile1_rxreset1_i                : std_logic;
    signal  tile1_rxbufreset1_i             : std_logic;

    signal  tile1_gtp0_cc_2b_1skp_cco_i     : std_logic_vector(6 downto 0);


    -- ground and tied_to_vcc_i signals
    signal  tied_to_ground_i                :   std_logic;
    signal  tied_to_ground_vec_i            :   std_logic_vector(63 downto 0);
    signal  tied_to_vcc_i                   :   std_logic;


--*************************** Component Declarations **************************

component ROCKETIO_WRAPPER_TILE
generic
(
    -- Simulation attributes
    TILE_SIM_MODE                : string    := "FAST"; -- Set to Fast Functional Simulation Model
    TILE_SIM_GTXRESET_SPEEDUP    : integer   := 0; -- Set to 1 to speed up sim reset
    TILE_SIM_PLL_PERDIV2         : bit_vector:= x"140"; -- Set to the VCO Unit Interval time

    -- Channel bonding attributes
    TILE_CHAN_BOND_MODE_0        : string    := "OFF";  -- "MASTER", "SLAVE", or "OFF"
    TILE_CHAN_BOND_LEVEL_0       : integer   := 0;     -- 0 to 7. See UG for details

    TILE_CHAN_BOND_MODE_1        : string    := "OFF";  -- "MASTER", "SLAVE", or "OFF"
    TILE_CHAN_BOND_LEVEL_1       : integer   := 0      -- 0 to 7. See UG for details
);
port
(
    ------------------------ Loopback and Powerdown Ports ----------------------
    LOOPBACK0_IN                            : in   std_logic_vector(2 downto 0);
    LOOPBACK1_IN                            : in   std_logic_vector(2 downto 0);
    RXPOWERDOWN0_IN                         : in   std_logic_vector(1 downto 0);
    RXPOWERDOWN1_IN                         : in   std_logic_vector(1 downto 0);
    TXPOWERDOWN0_IN                         : in   std_logic_vector(1 downto 0);
    TXPOWERDOWN1_IN                         : in   std_logic_vector(1 downto 0);
    ----------------------- Receive Ports - 8b10b Decoder ----------------------
    RXCHARISCOMMA0_OUT                      : out  std_logic_vector(1 downto 0);
    RXCHARISCOMMA1_OUT                      : out  std_logic_vector(1 downto 0);
    RXCHARISK0_OUT                          : out  std_logic_vector(1 downto 0);
    RXCHARISK1_OUT                          : out  std_logic_vector(1 downto 0);
    RXDISPERR0_OUT                          : out  std_logic_vector(1 downto 0);
    RXDISPERR1_OUT                          : out  std_logic_vector(1 downto 0);
    RXNOTINTABLE0_OUT                       : out  std_logic_vector(1 downto 0);
    RXNOTINTABLE1_OUT                       : out  std_logic_vector(1 downto 0);
    RXRUNDISP0_OUT                          : out  std_logic_vector(1 downto 0);
    RXRUNDISP1_OUT                          : out  std_logic_vector(1 downto 0);
    ------------------- Receive Ports - Channel Bonding Ports ------------------
    RXCHANBONDSEQ0_OUT                      : out  std_logic;
    RXCHANBONDSEQ1_OUT                      : out  std_logic;
    RXCHBONDI0_IN                           : in   std_logic_vector(3 downto 0);
    RXCHBONDI1_IN                           : in   std_logic_vector(3 downto 0);
    RXCHBONDO0_OUT                          : out  std_logic_vector(3 downto 0);
    RXCHBONDO1_OUT                          : out  std_logic_vector(3 downto 0);
    RXENCHANSYNC0_IN                        : in   std_logic;
    RXENCHANSYNC1_IN                        : in   std_logic;
    ------------------- Receive Ports - Clock Correction Ports -----------------
    RXCLKCORCNT0_OUT                        : out  std_logic_vector(2 downto 0);
    RXCLKCORCNT1_OUT                        : out  std_logic_vector(2 downto 0);
    --------------- Receive Ports - Comma Detection and Alignment --------------
    RXBYTEISALIGNED0_OUT                    : out  std_logic;
    RXBYTEISALIGNED1_OUT                    : out  std_logic;
    RXBYTEREALIGN0_OUT                      : out  std_logic;
    RXBYTEREALIGN1_OUT                      : out  std_logic;
    RXCOMMADET0_OUT                         : out  std_logic;
    RXCOMMADET1_OUT                         : out  std_logic;
    RXENMCOMMAALIGN0_IN                     : in   std_logic;
    RXENMCOMMAALIGN1_IN                     : in   std_logic;
    RXENPCOMMAALIGN0_IN                     : in   std_logic;
    RXENPCOMMAALIGN1_IN                     : in   std_logic;
    ------------------- Receive Ports - RX Data Path interface -----------------
    RXDATA0_OUT                             : out  std_logic_vector(15 downto 0);
    RXDATA1_OUT                             : out  std_logic_vector(15 downto 0);
    RXRECCLK0_OUT                           : out  std_logic;
    RXRECCLK1_OUT                           : out  std_logic;
    RXRESET0_IN                             : in   std_logic;
    RXRESET1_IN                             : in   std_logic;
    RXUSRCLK0_IN                            : in   std_logic;
    RXUSRCLK1_IN                            : in   std_logic;
    RXUSRCLK20_IN                           : in   std_logic;
    RXUSRCLK21_IN                           : in   std_logic;
    ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    RXCDRRESET0_IN                          : in   std_logic;
    RXCDRRESET1_IN                          : in   std_logic;
    RXELECIDLE0_OUT                         : out  std_logic;
    RXELECIDLE1_OUT                         : out  std_logic;
    RXN0_IN                                 : in   std_logic;
    RXN1_IN                                 : in   std_logic;
    RXP0_IN                                 : in   std_logic;
    RXP1_IN                                 : in   std_logic;
    -------- Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
    RXBUFRESET0_IN                          : in   std_logic;
    RXBUFRESET1_IN                          : in   std_logic;
    RXBUFSTATUS0_OUT                        : out  std_logic_vector(2 downto 0);
    RXBUFSTATUS1_OUT                        : out  std_logic_vector(2 downto 0);
    RXCHANISALIGNED0_OUT                    : out  std_logic;
    RXCHANISALIGNED1_OUT                    : out  std_logic;
    RXCHANREALIGN0_OUT                      : out  std_logic;
    RXCHANREALIGN1_OUT                      : out  std_logic;
    --------------- Receive Ports - RX Loss-of-sync State Machine --------------
    RXLOSSOFSYNC0_OUT                       : out  std_logic_vector(1 downto 0);
    RXLOSSOFSYNC1_OUT                       : out  std_logic_vector(1 downto 0);
    -------------- Receive Ports - RX Pipe Control for PCI Express -------------
    RXVALID0_OUT                            : out  std_logic;
    RXVALID1_OUT                            : out  std_logic;
    -------------- Receive Ports - polarity  -----------------------------------
    RXPOLARITY0                             : in   std_logic;
    RXPOLARITY1                             : in   std_logic;    
    ------------- Shared Ports - Dynamic Reconfiguration Port (DRP) ------------
    DADDR_IN                                : in   std_logic_vector(6 downto 0);
    DCLK_IN                                 : in   std_logic;
    DEN_IN                                  : in   std_logic;
    DI_IN                                   : in   std_logic_vector(15 downto 0);
    DO_OUT                                  : out  std_logic_vector(15 downto 0);
    DRDY_OUT                                : out  std_logic;
    DWE_IN                                  : in   std_logic;
    --------------------- Shared Ports - Tile and PLL Ports --------------------
    CLKIN_IN                                : in   std_logic;
    GTXRESET_IN                             : in   std_logic;
    PLLLKDET_OUT                            : out  std_logic;
    REFCLKOUT_OUT                           : out  std_logic;
    RESETDONE0_OUT                          : out  std_logic;
    RESETDONE1_OUT                          : out  std_logic;
    ---------------- Transmit Ports - 8b10b Encoder Control Ports --------------
    TXCHARISK0_IN                           : in   std_logic_vector(1 downto 0);
    TXCHARISK1_IN                           : in   std_logic_vector(1 downto 0);
    ------------------ Transmit Ports - TX Data Path interface -----------------
    TXDATA0_IN                              : in   std_logic_vector(15 downto 0);
    TXDATA1_IN                              : in   std_logic_vector(15 downto 0);
    TXRESET0_IN                             : in   std_logic;
    TXRESET1_IN                             : in   std_logic;
    TXUSRCLK0_IN                            : in   std_logic;
    TXUSRCLK1_IN                            : in   std_logic;
    TXUSRCLK20_IN                           : in   std_logic;
    TXUSRCLK21_IN                           : in   std_logic;
    --------------- Transmit Ports - TX Driver and OOB signalling --------------
    TXN0_OUT                                : out  std_logic;
    TXN1_OUT                                : out  std_logic;
    TXP0_OUT                                : out  std_logic;
    TXP1_OUT                                : out  std_logic;
    -------- Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
    TXENPMAPHASEALIGN0_IN                   : in   std_logic;
    TXENPMAPHASEALIGN1_IN                   : in   std_logic;
    TXPMASETPHASE0_IN                       : in   std_logic;
    TXPMASETPHASE1_IN                       : in   std_logic;
    -------------------- Transmit Ports - polarity  ----------------------------
    TXPOLARITY0                             : in   std_logic;
    TXPOLARITY1                             : in   std_logic;
    ----------------- Transmit Ports - TX Ports for PCI Express ----------------
    TXELECIDLE0_IN                          : in   std_logic;
    TXELECIDLE1_IN                          : in   std_logic


);
end component;

component CC_2B_1SKP
generic
(
    CC_CHAR                                 : in  std_logic_vector(7 downto 0) := X"1C";
    ALIGN_CHAR                              : in  std_logic_vector(7 downto 0) := X"7C";
    CHAN_BOND_MODE                          : in  string := "OFF";
    ALIGN_PARALLEL_CHECK                    : in  bit := '1';
    USE_AUTORECOVER                         : in  bit := '1';
    FIFO_ALMOST_EMPTY_OFFSET                : in  bit_vector := X"005";
    FIFO_ALMOST_FULL_OFFSET                 : in  bit_vector := X"1F2" --498
);
port
(
    GT_RXDATA                               : in   std_logic_vector(15 downto 0);
    GT_RXCHARISK                            : in   std_logic_vector(1  downto 0);
    GT_RXCHARISCOMMA                        : in   std_logic_vector(1  downto 0);
    GT_RXRUNDISP                            : in   std_logic_vector(1  downto 0);
    GT_RXNOTINTABLE                         : in   std_logic_vector(1  downto 0);
    GT_RXDISPERR                            : in   std_logic_vector(1  downto 0);
    GT_RXBUFSTATUS                          : in   std_logic_vector(2  downto 0);
    GT_RXCLKCORCNT                          : in   std_logic_vector(2  downto 0);
    GT_RXCHANBONDSEQ                        : in   std_logic;
    GT_RXCHANISALIGNED                      : in   std_logic;
    GT_RXCHANREALIGN                        : in   std_logic;
    GT_RXLOSSOFSYNC                         : in   std_logic_vector(1  downto 0);
    GT_RXVALID                              : in   std_logic;
    GT_RXUSRCLK2                            : in   std_logic;
    USER_RXUSRCLK2                          : in   std_logic;
    RESET                                   : in   std_logic;
    CCI                                     : in   std_logic_vector(6 downto 0);

    USER_RXDATA                             : out  std_logic_vector(15 downto 0);
    USER_RXCHARISK                          : out  std_logic_vector(1 downto 0);
    USER_RXCHARISCOMMA                      : out  std_logic_vector(1 downto 0);
    USER_RXRUNDISP                          : out  std_logic_vector(1 downto 0);
    USER_RXNOTINTABLE                       : out  std_logic_vector(1 downto 0);
    USER_RXDISPERR                          : out  std_logic_vector(1 downto 0);
    USER_RXBUFSTATUS                        : out  std_logic_vector(2 downto 0);
    USER_RXCLKCORCNT                        : out  std_logic_vector(2 downto 0);
    USER_RXCHANBONDSEQ                      : out  std_logic;
    USER_RXCHANISALIGNED                    : out  std_logic;
    USER_RXCHANREALIGN                      : out  std_logic;
    USER_RXLOSSOFSYNC                       : out  std_logic_vector(1 downto 0);
    USER_RXVALID                            : out  std_logic;
    CCO                                     : out  std_logic_vector(6 downto 0)
);
end component;


--********************************* Main Body of Code**************************

begin

    tied_to_ground_i                    <= '0';
    tied_to_ground_vec_i(63 downto 0)   <= (others => '0');
    tied_to_vcc_i                       <= '1';

    --------------------------- Tile Instances  -------------------------------

GEN_NO_SWAP0: if (not CH01_SWAP) generate
    --_________________________________________________________________________
    --_________________________________________________________________________
    --TILE0  (Location)

    tile0_rocketio_wrapper_i : ROCKETIO_WRAPPER_TILE
    generic map
    (
        -- Simulation attributes
        TILE_SIM_MODE                => WRAPPER_SIM_MODE,
        TILE_SIM_GTXRESET_SPEEDUP    => WRAPPER_SIM_GTXRESET_SPEEDUP,
        TILE_SIM_PLL_PERDIV2         => WRAPPER_SIM_PLL_PERDIV2,

        -- Channel bonding attributes
        TILE_CHAN_BOND_MODE_0        => "SLAVE",
        TILE_CHAN_BOND_LEVEL_0       => 0,

        TILE_CHAN_BOND_MODE_1        => "SLAVE",
        TILE_CHAN_BOND_LEVEL_1       => 0
    )
    port map
    (
        ------------------------ Loopback and Powerdown Ports ----------------------
        LOOPBACK0_IN                    =>      TILE0_LOOPBACK0_IN,
        LOOPBACK1_IN                    =>      TILE0_LOOPBACK1_IN,
        RXPOWERDOWN0_IN                 =>      TILE0_RXPOWERDOWN0_IN,
        RXPOWERDOWN1_IN                 =>      TILE0_RXPOWERDOWN1_IN,
        TXPOWERDOWN0_IN                 =>      TILE0_TXPOWERDOWN0_IN,
        TXPOWERDOWN1_IN                 =>      TILE0_TXPOWERDOWN1_IN,
        ----------------------- Receive Ports - 8b10b Decoder ----------------------
        RXCHARISCOMMA0_OUT              =>      tile0_rxchariscomma0_i,
        RXCHARISCOMMA1_OUT              =>      tile0_rxchariscomma1_i,
        RXCHARISK0_OUT                  =>      tile0_rxcharisk0_i,
        RXCHARISK1_OUT                  =>      tile0_rxcharisk1_i,
        RXDISPERR0_OUT                  =>      tile0_rxdisperr0_i,
        RXDISPERR1_OUT                  =>      tile0_rxdisperr1_i,
        RXNOTINTABLE0_OUT               =>      tile0_rxnotintable0_i,
        RXNOTINTABLE1_OUT               =>      tile0_rxnotintable1_i,
        RXRUNDISP0_OUT                  =>      tile0_rxrundisp0_i,
        RXRUNDISP1_OUT                  =>      tile0_rxrundisp1_i,
        ------------------- Receive Ports - Channel Bonding Ports ------------------
        RXCHANBONDSEQ0_OUT              =>      tile0_rxchanbondseq0_i,
        RXCHANBONDSEQ1_OUT              =>      tile0_rxchanbondseq1_i,
        RXCHBONDI0_IN                   =>      tile1_rxchbondo1_i,
        RXCHBONDI1_IN                   =>      tile1_rxchbondo1_i,
        RXCHBONDO0_OUT                  =>      tile0_rxchbondo0_i,
        RXCHBONDO1_OUT                  =>      tile0_rxchbondo1_i,
        RXENCHANSYNC0_IN                =>      TILE0_RXENCHANSYNC0_IN,
        RXENCHANSYNC1_IN                =>      TILE0_RXENCHANSYNC1_IN,
        ------------------- Receive Ports - Clock Correction Ports -----------------
        RXCLKCORCNT0_OUT                =>      tile0_rxclkcorcnt0_i,
        RXCLKCORCNT1_OUT                =>      tile0_rxclkcorcnt1_i,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        RXBYTEISALIGNED0_OUT            =>      TILE0_RXBYTEISALIGNED0_OUT,
        RXBYTEISALIGNED1_OUT            =>      TILE0_RXBYTEISALIGNED1_OUT,
        RXBYTEREALIGN0_OUT              =>      TILE0_RXBYTEREALIGN0_OUT,
        RXBYTEREALIGN1_OUT              =>      TILE0_RXBYTEREALIGN1_OUT,
        RXCOMMADET0_OUT                 =>      TILE0_RXCOMMADET0_OUT,
        RXCOMMADET1_OUT                 =>      TILE0_RXCOMMADET1_OUT,
        RXENMCOMMAALIGN0_IN             =>      TILE0_RXENMCOMMAALIGN0_IN,
        RXENMCOMMAALIGN1_IN             =>      TILE0_RXENMCOMMAALIGN1_IN,
        RXENPCOMMAALIGN0_IN             =>      TILE0_RXENPCOMMAALIGN0_IN,
        RXENPCOMMAALIGN1_IN             =>      TILE0_RXENPCOMMAALIGN1_IN,
        ------------------- Receive Ports - RX Data Path interface -----------------
        RXDATA0_OUT                     =>      tile0_rxdata0_i,
        RXDATA1_OUT                     =>      tile0_rxdata1_i,
        RXRECCLK0_OUT                   =>      tile0_rxrecclk0_i,
        RXRECCLK1_OUT                   =>      tile0_rxrecclk1_i,
        RXRESET0_IN                     =>      tile0_rxreset0_i,
        RXRESET1_IN                     =>      tile0_rxreset1_i,
        RXUSRCLK0_IN                    =>      tile1_rxrecclk0_bufg_i,
        RXUSRCLK1_IN                    =>      tile1_rxrecclk0_bufg_i,
        RXUSRCLK20_IN                   =>      tile1_rxrecclk0_bufg_i,
        RXUSRCLK21_IN                   =>      tile1_rxrecclk0_bufg_i,
        ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        RXCDRRESET0_IN                  =>      TILE0_RXCDRRESET0_IN,
        RXCDRRESET1_IN                  =>      TILE0_RXCDRRESET1_IN,
        RXELECIDLE0_OUT                 =>      TILE0_RXELECIDLE0_OUT,
        RXELECIDLE1_OUT                 =>      TILE0_RXELECIDLE1_OUT,
        RXN0_IN                         =>      TILE0_RXN0_IN,
        RXN1_IN                         =>      TILE0_RXN1_IN,
        RXP0_IN                         =>      TILE0_RXP0_IN,
        RXP1_IN                         =>      TILE0_RXP1_IN,
        -------- Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
        RXBUFRESET0_IN                  =>      tile0_rxbufreset0_i,
        RXBUFRESET1_IN                  =>      tile0_rxbufreset1_i,
        RXBUFSTATUS0_OUT                =>      tile0_rxbufstatus0_i,
        RXBUFSTATUS1_OUT                =>      tile0_rxbufstatus1_i,
        RXCHANISALIGNED0_OUT            =>      tile0_rxchanisaligned0_i,
        RXCHANISALIGNED1_OUT            =>      tile0_rxchanisaligned1_i,
        RXCHANREALIGN0_OUT              =>      tile0_rxchanrealign0_i,
        RXCHANREALIGN1_OUT              =>      tile0_rxchanrealign1_i,
        --------------- Receive Ports - RX Loss-of-sync State Machine --------------
        RXLOSSOFSYNC0_OUT               =>      tile0_rxlossofsync0_i,
        RXLOSSOFSYNC1_OUT               =>      tile0_rxlossofsync1_i,
        -------------- Receive Ports - polarity  -----------------------------------
        RXPOLARITY0                     =>      TILE0_RXPOLARITY0,
        RXPOLARITY1                     =>      TILE0_RXPOLARITY1,    
        -------------- Receive Ports - RX Pipe Control for PCI Express -------------
        RXVALID0_OUT                    =>      tile0_rxvalid0_i,
        RXVALID1_OUT                    =>      tile0_rxvalid1_i,
        ------------- Shared Ports - Dynamic Reconfiguration Port (DRP) ------------
        DADDR_IN                        =>      TILE0_DADDR_IN,
        DCLK_IN                         =>      TILE0_DCLK_IN,
        DEN_IN                          =>      TILE0_DEN_IN,
        DI_IN                           =>      TILE0_DI_IN,
        DO_OUT                          =>      TILE0_DO_OUT,
        DRDY_OUT                        =>      TILE0_DRDY_OUT,
        DWE_IN                          =>      TILE0_DWE_IN,
        --------------------- Shared Ports - Tile and PLL Ports --------------------
        CLKIN_IN                        =>      TILE0_CLKIN_IN,
        GTXRESET_IN                     =>      TILE0_GTXRESET_IN,
        PLLLKDET_OUT                    =>      TILE0_PLLLKDET_OUT,
        REFCLKOUT_OUT                   =>      TILE0_REFCLKOUT_OUT,
        RESETDONE0_OUT                  =>      tile0_resetdone0_i,
        RESETDONE1_OUT                  =>      tile0_resetdone1_i,
        ---------------- Transmit Ports - 8b10b Encoder Control Ports --------------
        TXCHARISK0_IN                   =>      TILE0_TXCHARISK0_IN,
        TXCHARISK1_IN                   =>      TILE0_TXCHARISK1_IN,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        TXDATA0_IN                      =>      TILE0_TXDATA0_IN,
        TXDATA1_IN                      =>      TILE0_TXDATA1_IN,
        TXRESET0_IN                     =>      TILE0_TXRESET0_IN,
        TXRESET1_IN                     =>      TILE0_TXRESET1_IN,
        TXUSRCLK0_IN                    =>      TILE0_TXUSRCLK0_IN,
        TXUSRCLK1_IN                    =>      TILE0_TXUSRCLK1_IN,
        TXUSRCLK20_IN                   =>      TILE0_TXUSRCLK20_IN,
        TXUSRCLK21_IN                   =>      TILE0_TXUSRCLK21_IN,
        --------------- Transmit Ports - TX Driver and OOB signalling --------------
        TXN0_OUT                        =>      TILE0_TXN0_OUT,
        TXN1_OUT                        =>      TILE0_TXN1_OUT,
        TXP0_OUT                        =>      TILE0_TXP0_OUT,
        TXP1_OUT                        =>      TILE0_TXP1_OUT,
        -------- Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
        TXENPMAPHASEALIGN0_IN           =>      TILE0_TXENPMAPHASEALIGN0_IN,
        TXENPMAPHASEALIGN1_IN           =>      TILE0_TXENPMAPHASEALIGN1_IN,
        TXPMASETPHASE0_IN               =>      TILE0_TXPMASETPHASE0_IN,
        TXPMASETPHASE1_IN               =>      TILE0_TXPMASETPHASE1_IN,
        -------------------- Transmit Ports - polarity  ----------------------------
        TXPOLARITY0                     =>      TILE0_TXPOLARITY0,
        TXPOLARITY1                     =>      TILE0_TXPOLARITY1,
        ----------------- Transmit Ports - TX Ports for PCI Express ----------------
        TXELECIDLE0_IN                  =>      TILE0_TXELECIDLE0_IN,
        TXELECIDLE1_IN                  =>      TILE0_TXELECIDLE1_IN

    );
end generate;

GEN_SWAP0: if (CH01_SWAP) generate
    --_________________________________________________________________________
    --_________________________________________________________________________
    --TILE0  (Location)
    tile0_rocketio_wrapper_i : ROCKETIO_WRAPPER_TILE
    generic map
    (
        -- Simulation attributes
        TILE_SIM_MODE                => WRAPPER_SIM_MODE,
        TILE_SIM_GTXRESET_SPEEDUP    => WRAPPER_SIM_GTXRESET_SPEEDUP,
        TILE_SIM_PLL_PERDIV2         => WRAPPER_SIM_PLL_PERDIV2,

        -- Channel bonding attributes
        TILE_CHAN_BOND_MODE_0        => "SLAVE",
        TILE_CHAN_BOND_LEVEL_0       => 0,

        TILE_CHAN_BOND_MODE_1        => "SLAVE",
        TILE_CHAN_BOND_LEVEL_1       => 0
    )
    port map
    (
        ------------------------ Loopback and Powerdown Ports ----------------------
        LOOPBACK0_IN                    =>      TILE0_LOOPBACK1_IN,
        LOOPBACK1_IN                    =>      TILE0_LOOPBACK0_IN,
        RXPOWERDOWN0_IN                 =>      TILE0_RXPOWERDOWN1_IN,
        RXPOWERDOWN1_IN                 =>      TILE0_RXPOWERDOWN0_IN,
        TXPOWERDOWN0_IN                 =>      TILE0_TXPOWERDOWN1_IN,
        TXPOWERDOWN1_IN                 =>      TILE0_TXPOWERDOWN0_IN,
        ----------------------- Receive Ports - 8b10b Decoder ----------------------
        RXCHARISCOMMA0_OUT              =>      tile0_rxchariscomma1_i,
        RXCHARISCOMMA1_OUT              =>      tile0_rxchariscomma0_i,
        RXCHARISK0_OUT                  =>      tile0_rxcharisk1_i,
        RXCHARISK1_OUT                  =>      tile0_rxcharisk0_i,
        RXDISPERR0_OUT                  =>      tile0_rxdisperr1_i,
        RXDISPERR1_OUT                  =>      tile0_rxdisperr0_i,
        RXNOTINTABLE0_OUT               =>      tile0_rxnotintable1_i,
        RXNOTINTABLE1_OUT               =>      tile0_rxnotintable0_i,
        RXRUNDISP0_OUT                  =>      tile0_rxrundisp1_i,
        RXRUNDISP1_OUT                  =>      tile0_rxrundisp0_i,
        ------------------- Receive Ports - Channel Bonding Ports ------------------
        RXCHANBONDSEQ0_OUT              =>      tile0_rxchanbondseq1_i,
        RXCHANBONDSEQ1_OUT              =>      tile0_rxchanbondseq0_i,
        RXCHBONDI0_IN                   =>      tile1_rxchbondo1_i,
        RXCHBONDI1_IN                   =>      tile1_rxchbondo1_i,
        RXCHBONDO0_OUT                  =>      tile0_rxchbondo1_i,
        RXCHBONDO1_OUT                  =>      tile0_rxchbondo0_i,
        RXENCHANSYNC0_IN                =>      TILE0_RXENCHANSYNC1_IN,
        RXENCHANSYNC1_IN                =>      TILE0_RXENCHANSYNC0_IN,
        ------------------- Receive Ports - Clock Correction Ports -----------------
        RXCLKCORCNT0_OUT                =>      tile0_rxclkcorcnt1_i,
        RXCLKCORCNT1_OUT                =>      tile0_rxclkcorcnt0_i,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        RXBYTEISALIGNED0_OUT            =>      TILE0_RXBYTEISALIGNED1_OUT,
        RXBYTEISALIGNED1_OUT            =>      TILE0_RXBYTEISALIGNED0_OUT,
        RXBYTEREALIGN0_OUT              =>      TILE0_RXBYTEREALIGN1_OUT,
        RXBYTEREALIGN1_OUT              =>      TILE0_RXBYTEREALIGN0_OUT,
        RXCOMMADET0_OUT                 =>      TILE0_RXCOMMADET1_OUT,
        RXCOMMADET1_OUT                 =>      TILE0_RXCOMMADET0_OUT,
        RXENMCOMMAALIGN0_IN             =>      TILE0_RXENMCOMMAALIGN1_IN,
        RXENMCOMMAALIGN1_IN             =>      TILE0_RXENMCOMMAALIGN0_IN,
        RXENPCOMMAALIGN0_IN             =>      TILE0_RXENPCOMMAALIGN1_IN,
        RXENPCOMMAALIGN1_IN             =>      TILE0_RXENPCOMMAALIGN0_IN,
        ------------------- Receive Ports - RX Data Path interface -----------------
        RXDATA0_OUT                     =>      tile0_rxdata1_i,
        RXDATA1_OUT                     =>      tile0_rxdata0_i,
        RXRECCLK0_OUT                   =>      tile0_rxrecclk1_i,
        RXRECCLK1_OUT                   =>      tile0_rxrecclk0_i,
        RXRESET0_IN                     =>      tile0_rxreset1_i,
        RXRESET1_IN                     =>      tile0_rxreset0_i,
        RXUSRCLK0_IN                    =>      tile1_rxrecclk0_bufg_i,
        RXUSRCLK1_IN                    =>      tile1_rxrecclk0_bufg_i,
        RXUSRCLK20_IN                   =>      tile1_rxrecclk0_bufg_i,
        RXUSRCLK21_IN                   =>      tile1_rxrecclk0_bufg_i,
        ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        RXCDRRESET0_IN                  =>      TILE0_RXCDRRESET1_IN,
        RXCDRRESET1_IN                  =>      TILE0_RXCDRRESET0_IN,
        RXELECIDLE0_OUT                 =>      TILE0_RXELECIDLE1_OUT,
        RXELECIDLE1_OUT                 =>      TILE0_RXELECIDLE0_OUT,
        RXN0_IN                         =>      TILE0_RXN1_IN,
        RXN1_IN                         =>      TILE0_RXN0_IN,
        RXP0_IN                         =>      TILE0_RXP1_IN,
        RXP1_IN                         =>      TILE0_RXP0_IN,
        -------- Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
        RXBUFRESET0_IN                  =>      tile0_rxbufreset1_i,
        RXBUFRESET1_IN                  =>      tile0_rxbufreset0_i,
        RXBUFSTATUS0_OUT                =>      tile0_rxbufstatus1_i,
        RXBUFSTATUS1_OUT                =>      tile0_rxbufstatus0_i,
        RXCHANISALIGNED0_OUT            =>      tile0_rxchanisaligned1_i,
        RXCHANISALIGNED1_OUT            =>      tile0_rxchanisaligned0_i,
        RXCHANREALIGN0_OUT              =>      tile0_rxchanrealign1_i,
        RXCHANREALIGN1_OUT              =>      tile0_rxchanrealign0_i,
        --------------- Receive Ports - RX Loss-of-sync State Machine --------------
        RXLOSSOFSYNC0_OUT               =>      tile0_rxlossofsync1_i,
        RXLOSSOFSYNC1_OUT               =>      tile0_rxlossofsync0_i,
        -------------- Receive Ports - polarity  -----------------------------------
        RXPOLARITY0                     =>      TILE0_RXPOLARITY1,
        RXPOLARITY1                     =>      TILE0_RXPOLARITY0,            
        -------------- Receive Ports - RX Pipe Control for PCI Express -------------
        RXVALID0_OUT                    =>      tile0_rxvalid1_i,
        RXVALID1_OUT                    =>      tile0_rxvalid0_i,
        ------------- Shared Ports - Dynamic Reconfiguration Port (DRP) ------------
        DADDR_IN                        =>      TILE0_DADDR_IN,
        DCLK_IN                         =>      TILE0_DCLK_IN,
        DEN_IN                          =>      TILE0_DEN_IN,
        DI_IN                           =>      TILE0_DI_IN,
        DO_OUT                          =>      TILE0_DO_OUT,
        DRDY_OUT                        =>      TILE0_DRDY_OUT,
        DWE_IN                          =>      TILE0_DWE_IN,
        --------------------- Shared Ports - Tile and PLL Ports --------------------
        CLKIN_IN                        =>      TILE0_CLKIN_IN,
        GTXRESET_IN                     =>      TILE0_GTXRESET_IN,
        PLLLKDET_OUT                    =>      TILE0_PLLLKDET_OUT,
        REFCLKOUT_OUT                   =>      TILE0_REFCLKOUT_OUT,
        RESETDONE0_OUT                  =>      tile0_resetdone1_i,
        RESETDONE1_OUT                  =>      tile0_resetdone0_i,
        ---------------- Transmit Ports - 8b10b Encoder Control Ports --------------
        TXCHARISK0_IN                   =>      TILE0_TXCHARISK1_IN,
        TXCHARISK1_IN                   =>      TILE0_TXCHARISK0_IN,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        TXDATA0_IN                      =>      TILE0_TXDATA1_IN,
        TXDATA1_IN                      =>      TILE0_TXDATA0_IN,
        TXRESET0_IN                     =>      TILE0_TXRESET1_IN,
        TXRESET1_IN                     =>      TILE0_TXRESET0_IN,
        TXUSRCLK0_IN                    =>      TILE0_TXUSRCLK1_IN,
        TXUSRCLK1_IN                    =>      TILE0_TXUSRCLK0_IN,
        TXUSRCLK20_IN                   =>      TILE0_TXUSRCLK21_IN,
        TXUSRCLK21_IN                   =>      TILE0_TXUSRCLK20_IN,
        --------------- Transmit Ports - TX Driver and OOB signalling --------------
        TXN0_OUT                        =>      TILE0_TXN1_OUT,
        TXN1_OUT                        =>      TILE0_TXN0_OUT,
        TXP0_OUT                        =>      TILE0_TXP1_OUT,
        TXP1_OUT                        =>      TILE0_TXP0_OUT,
        -------- Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
        TXENPMAPHASEALIGN0_IN           =>      TILE0_TXENPMAPHASEALIGN1_IN,
        TXENPMAPHASEALIGN1_IN           =>      TILE0_TXENPMAPHASEALIGN0_IN,
        TXPMASETPHASE0_IN               =>      TILE0_TXPMASETPHASE1_IN,
        TXPMASETPHASE1_IN               =>      TILE0_TXPMASETPHASE0_IN,
        -------------------- Transmit Ports - polarity  ----------------------------
        TXPOLARITY0                     =>      TILE0_TXPOLARITY1,
        TXPOLARITY1                     =>      TILE0_TXPOLARITY0,
        ----------------- Transmit Ports - TX Ports for PCI Express ----------------
        TXELECIDLE0_IN                  =>      TILE0_TXELECIDLE1_IN,
        TXELECIDLE1_IN                  =>      TILE0_TXELECIDLE0_IN

    );
end generate;

    --_________________________________________________________________________
    --_________________________________________________________________________
    --TILE0 GTP0
    tile0_gtp0_cc_2b_1skp_i : CC_2B_1SKP
    generic map
    (
        CC_CHAR                      => x"1c",
        ALIGN_CHAR                   => x"7c",
        CHAN_BOND_MODE               => "SLAVE",
        ALIGN_PARALLEL_CHECK         => '1'
    )
    port map
    (
        -- Write Interface on the RXRECCLK
        GT_RXDATA                       =>      tile0_rxdata0_i,
        GT_RXCHARISK                    =>      tile0_rxcharisk0_i,
        GT_RXCHARISCOMMA                =>      tile0_rxchariscomma0_i,
        GT_RXRUNDISP                    =>      tile0_rxrundisp0_i,
        GT_RXNOTINTABLE                 =>      tile0_rxnotintable0_i,
        GT_RXDISPERR                    =>      tile0_rxdisperr0_i,
        GT_RXBUFSTATUS                  =>      tile0_rxbufstatus0_i,
        GT_RXCLKCORCNT                  =>      tile0_rxclkcorcnt0_i,
        GT_RXCHANBONDSEQ                =>      tile0_rxchanbondseq0_i,
        GT_RXCHANISALIGNED              =>      tile0_rxchanisaligned0_i,
        GT_RXCHANREALIGN                =>      tile0_rxchanrealign0_i,
        GT_RXLOSSOFSYNC                 =>      tile0_rxlossofsync0_i,
        GT_RXVALID                      =>      tile0_rxvalid0_i,
        GT_RXUSRCLK2                    =>      tile1_rxrecclk0_bufg_i,

        -- Read Interface on the RXUSRCLK2
        USER_RXDATA                     =>      TILE0_RXDATA0_OUT,
        USER_RXCHARISK                  =>      TILE0_RXCHARISK0_OUT,
        USER_RXCHARISCOMMA              =>      TILE0_RXCHARISCOMMA0_OUT,
        USER_RXRUNDISP                  =>      open,
        USER_RXNOTINTABLE               =>      TILE0_RXNOTINTABLE0_OUT,
        USER_RXDISPERR                  =>      TILE0_RXDISPERR0_OUT,
        USER_RXBUFSTATUS                =>      TILE0_RXBUFSTATUS0_OUT,
        USER_RXCLKCORCNT                =>      TILE0_RXCLKCORCNT0_OUT,
        USER_RXCHANBONDSEQ              =>      TILE0_RXCHANBONDSEQ0_OUT,
        USER_RXCHANISALIGNED            =>      TILE0_RXCHANISALIGNED0_OUT,
        USER_RXCHANREALIGN              =>      TILE0_RXCHANREALIGN0_OUT,
        USER_RXLOSSOFSYNC               =>      TILE0_RXLOSSOFSYNC0_OUT,
        USER_RXVALID                    =>      open,
        USER_RXUSRCLK2                  =>      TILE0_RXUSRCLK20_IN,

        -- Status and reset signals
        RESET                           =>      tied_to_ground_i,
        CCI                             =>      tile1_gtp0_cc_2b_1skp_cco_i,
        CCO                             =>      open
    );

    TILE0_RESETDONE0_OUT <= tile0_resetdone0_i;
    tile0_rxreset0_i <= TILE0_RXRESET0_IN;
    tile0_rxbufreset0_i <= TILE0_RXBUFRESET0_IN;
    
    --_________________________________________________________________________
    --_________________________________________________________________________
    --TILE0 GTP1
    tile0_gtp1_cc_2b_1skp_i : CC_2B_1SKP
    generic map
    (
        CC_CHAR                      => x"1c",
        ALIGN_CHAR                   => x"7c",
        CHAN_BOND_MODE               => "SLAVE",
        ALIGN_PARALLEL_CHECK         => '1'
    )
    port map
    (
        -- Write Interface on the RXRECCLK
        GT_RXDATA                       =>      tile0_rxdata1_i,
        GT_RXCHARISK                    =>      tile0_rxcharisk1_i,
        GT_RXCHARISCOMMA                =>      tile0_rxchariscomma1_i,
        GT_RXRUNDISP                    =>      tile0_rxrundisp1_i,
        GT_RXNOTINTABLE                 =>      tile0_rxnotintable1_i,
        GT_RXDISPERR                    =>      tile0_rxdisperr1_i,
        GT_RXBUFSTATUS                  =>      tile0_rxbufstatus1_i,
        GT_RXCLKCORCNT                  =>      tile0_rxclkcorcnt1_i,
        GT_RXCHANBONDSEQ                =>      tile0_rxchanbondseq1_i,
        GT_RXCHANISALIGNED              =>      tile0_rxchanisaligned1_i,
        GT_RXCHANREALIGN                =>      tile0_rxchanrealign1_i,
        GT_RXLOSSOFSYNC                 =>      tile0_rxlossofsync1_i,
        GT_RXVALID                      =>      tile0_rxvalid1_i,
        GT_RXUSRCLK2                    =>      tile1_rxrecclk0_bufg_i,

        -- Read Interface on the RXUSRCLK2
        USER_RXDATA                     =>      TILE0_RXDATA1_OUT,
        USER_RXCHARISK                  =>      TILE0_RXCHARISK1_OUT,
        USER_RXCHARISCOMMA              =>      TILE0_RXCHARISCOMMA1_OUT,
        USER_RXRUNDISP                  =>      open,
        USER_RXNOTINTABLE               =>      TILE0_RXNOTINTABLE1_OUT,
        USER_RXDISPERR                  =>      TILE0_RXDISPERR1_OUT,
        USER_RXBUFSTATUS                =>      TILE0_RXBUFSTATUS1_OUT,
        USER_RXCLKCORCNT                =>      TILE0_RXCLKCORCNT1_OUT,
        USER_RXCHANBONDSEQ              =>      TILE0_RXCHANBONDSEQ1_OUT,
        USER_RXCHANISALIGNED            =>      TILE0_RXCHANISALIGNED1_OUT,
        USER_RXCHANREALIGN              =>      TILE0_RXCHANREALIGN1_OUT,
        USER_RXLOSSOFSYNC               =>      TILE0_RXLOSSOFSYNC1_OUT,
        USER_RXVALID                    =>      open,
        USER_RXUSRCLK2                  =>      TILE0_RXUSRCLK21_IN,

        -- Status and reset signals
        RESET                           =>      tied_to_ground_i,
        CCI                             =>      tile1_gtp0_cc_2b_1skp_cco_i,
        CCO                             =>      open
    );

    TILE0_RESETDONE1_OUT <= tile0_resetdone1_i;
    tile0_rxreset1_i <= TILE0_RXRESET1_IN;
    tile0_rxbufreset1_i <= TILE0_RXBUFRESET1_IN;

GEN_NO_SWAP1: if (not CH23_SWAP) generate
    --_________________________________________________________________________
    --_________________________________________________________________________
    --TILE1  (Location)

    tile1_rocketio_wrapper_i : ROCKETIO_WRAPPER_TILE
    generic map
    (
        -- Simulation attributes
        TILE_SIM_MODE                => WRAPPER_SIM_MODE,
        TILE_SIM_GTXRESET_SPEEDUP    => WRAPPER_SIM_GTXRESET_SPEEDUP,
        TILE_SIM_PLL_PERDIV2         => WRAPPER_SIM_PLL_PERDIV2,

        -- Channel bonding attributes
        TILE_CHAN_BOND_MODE_0        => "MASTER",
        TILE_CHAN_BOND_LEVEL_0       => 2,

        TILE_CHAN_BOND_MODE_1        => "SLAVE",
        TILE_CHAN_BOND_LEVEL_1       => 1
    )
    port map
    (
        ------------------------ Loopback and Powerdown Ports ----------------------
        LOOPBACK0_IN                    =>      TILE1_LOOPBACK0_IN,
        LOOPBACK1_IN                    =>      TILE1_LOOPBACK1_IN,
        RXPOWERDOWN0_IN                 =>      TILE1_RXPOWERDOWN0_IN,
        RXPOWERDOWN1_IN                 =>      TILE1_RXPOWERDOWN1_IN,
        TXPOWERDOWN0_IN                 =>      TILE1_TXPOWERDOWN0_IN,
        TXPOWERDOWN1_IN                 =>      TILE1_TXPOWERDOWN1_IN,
        ----------------------- Receive Ports - 8b10b Decoder ----------------------
        RXCHARISCOMMA0_OUT              =>      tile1_rxchariscomma0_i,
        RXCHARISCOMMA1_OUT              =>      tile1_rxchariscomma1_i,
        RXCHARISK0_OUT                  =>      tile1_rxcharisk0_i,
        RXCHARISK1_OUT                  =>      tile1_rxcharisk1_i,
        RXDISPERR0_OUT                  =>      tile1_rxdisperr0_i,
        RXDISPERR1_OUT                  =>      tile1_rxdisperr1_i,
        RXNOTINTABLE0_OUT               =>      tile1_rxnotintable0_i,
        RXNOTINTABLE1_OUT               =>      tile1_rxnotintable1_i,
        RXRUNDISP0_OUT                  =>      tile1_rxrundisp0_i,
        RXRUNDISP1_OUT                  =>      tile1_rxrundisp1_i,
        ------------------- Receive Ports - Channel Bonding Ports ------------------
        RXCHANBONDSEQ0_OUT              =>      tile1_rxchanbondseq0_i,
        RXCHANBONDSEQ1_OUT              =>      tile1_rxchanbondseq1_i,
        RXCHBONDI0_IN                   =>      tied_to_ground_vec_i(3 downto 0),
        RXCHBONDI1_IN                   =>      tile1_rxchbondo0_i,
        RXCHBONDO0_OUT                  =>      tile1_rxchbondo0_i,
        RXCHBONDO1_OUT                  =>      tile1_rxchbondo1_i,
        RXENCHANSYNC0_IN                =>      TILE1_RXENCHANSYNC0_IN,
        RXENCHANSYNC1_IN                =>      TILE1_RXENCHANSYNC1_IN,
        ------------------- Receive Ports - Clock Correction Ports -----------------
        RXCLKCORCNT0_OUT                =>      tile1_rxclkcorcnt0_i,
        RXCLKCORCNT1_OUT                =>      tile1_rxclkcorcnt1_i,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        RXBYTEISALIGNED0_OUT            =>      TILE1_RXBYTEISALIGNED0_OUT,
        RXBYTEISALIGNED1_OUT            =>      TILE1_RXBYTEISALIGNED1_OUT,
        RXBYTEREALIGN0_OUT              =>      TILE1_RXBYTEREALIGN0_OUT,
        RXBYTEREALIGN1_OUT              =>      TILE1_RXBYTEREALIGN1_OUT,
        RXCOMMADET0_OUT                 =>      TILE1_RXCOMMADET0_OUT,
        RXCOMMADET1_OUT                 =>      TILE1_RXCOMMADET1_OUT,
        RXENMCOMMAALIGN0_IN             =>      TILE1_RXENMCOMMAALIGN0_IN,
        RXENMCOMMAALIGN1_IN             =>      TILE1_RXENMCOMMAALIGN1_IN,
        RXENPCOMMAALIGN0_IN             =>      TILE1_RXENPCOMMAALIGN0_IN,
        RXENPCOMMAALIGN1_IN             =>      TILE1_RXENPCOMMAALIGN1_IN,
        ------------------- Receive Ports - RX Data Path interface -----------------
        RXDATA0_OUT                     =>      tile1_rxdata0_i,
        RXDATA1_OUT                     =>      tile1_rxdata1_i,
        RXRECCLK0_OUT                   =>      tile1_rxrecclk0_i,
        RXRECCLK1_OUT                   =>      tile1_rxrecclk1_i,
        RXRESET0_IN                     =>      tile1_rxreset0_i,
        RXRESET1_IN                     =>      tile1_rxreset1_i,
        RXUSRCLK0_IN                    =>      tile1_rxrecclk0_bufg_i,
        RXUSRCLK1_IN                    =>      tile1_rxrecclk0_bufg_i,
        RXUSRCLK20_IN                   =>      tile1_rxrecclk0_bufg_i,
        RXUSRCLK21_IN                   =>      tile1_rxrecclk0_bufg_i,
        ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        RXCDRRESET0_IN                  =>      TILE1_RXCDRRESET0_IN,
        RXCDRRESET1_IN                  =>      TILE1_RXCDRRESET1_IN,
        RXELECIDLE0_OUT                 =>      TILE1_RXELECIDLE0_OUT,
        RXELECIDLE1_OUT                 =>      TILE1_RXELECIDLE1_OUT,
        RXN0_IN                         =>      TILE1_RXN0_IN,
        RXN1_IN                         =>      TILE1_RXN1_IN,
        RXP0_IN                         =>      TILE1_RXP0_IN,
        RXP1_IN                         =>      TILE1_RXP1_IN,
        -------- Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
        RXBUFRESET0_IN                  =>      tile1_rxbufreset0_i,
        RXBUFRESET1_IN                  =>      tile1_rxbufreset1_i,
        RXBUFSTATUS0_OUT                =>      tile1_rxbufstatus0_i,
        RXBUFSTATUS1_OUT                =>      tile1_rxbufstatus1_i,
        RXCHANISALIGNED0_OUT            =>      tile1_rxchanisaligned0_i,
        RXCHANISALIGNED1_OUT            =>      tile1_rxchanisaligned1_i,
        RXCHANREALIGN0_OUT              =>      tile1_rxchanrealign0_i,
        RXCHANREALIGN1_OUT              =>      tile1_rxchanrealign1_i,
        --------------- Receive Ports - RX Loss-of-sync State Machine --------------
        RXLOSSOFSYNC0_OUT               =>      tile1_rxlossofsync0_i,
        RXLOSSOFSYNC1_OUT               =>      tile1_rxlossofsync1_i,
        -------------- Receive Ports - polarity  -----------------------------------
        RXPOLARITY0                     =>      TILE1_RXPOLARITY0,
        RXPOLARITY1                     =>      TILE1_RXPOLARITY1,
        -------------- Receive Ports - RX Pipe Control for PCI Express -------------
        RXVALID0_OUT                    =>      tile1_rxvalid0_i,
        RXVALID1_OUT                    =>      tile1_rxvalid1_i,
        ------------- Shared Ports - Dynamic Reconfiguration Port (DRP) ------------
        DADDR_IN                        =>      TILE1_DADDR_IN,
        DCLK_IN                         =>      TILE1_DCLK_IN,
        DEN_IN                          =>      TILE1_DEN_IN,
        DI_IN                           =>      TILE1_DI_IN,
        DO_OUT                          =>      TILE1_DO_OUT,
        DRDY_OUT                        =>      TILE1_DRDY_OUT,
        DWE_IN                          =>      TILE1_DWE_IN,
        --------------------- Shared Ports - Tile and PLL Ports --------------------
        CLKIN_IN                        =>      TILE1_CLKIN_IN,
        GTXRESET_IN                     =>      TILE1_GTXRESET_IN,
        PLLLKDET_OUT                    =>      TILE1_PLLLKDET_OUT,
        REFCLKOUT_OUT                   =>      TILE1_REFCLKOUT_OUT,
        RESETDONE0_OUT                  =>      tile1_resetdone0_i,
        RESETDONE1_OUT                  =>      tile1_resetdone1_i,
        ---------------- Transmit Ports - 8b10b Encoder Control Ports --------------
        TXCHARISK0_IN                   =>      TILE1_TXCHARISK0_IN,
        TXCHARISK1_IN                   =>      TILE1_TXCHARISK1_IN,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        TXDATA0_IN                      =>      TILE1_TXDATA0_IN,
        TXDATA1_IN                      =>      TILE1_TXDATA1_IN,
        TXRESET0_IN                     =>      TILE1_TXRESET0_IN,
        TXRESET1_IN                     =>      TILE1_TXRESET1_IN,
        TXUSRCLK0_IN                    =>      TILE1_TXUSRCLK0_IN,
        TXUSRCLK1_IN                    =>      TILE1_TXUSRCLK1_IN,
        TXUSRCLK20_IN                   =>      TILE1_TXUSRCLK20_IN,
        TXUSRCLK21_IN                   =>      TILE1_TXUSRCLK21_IN,
        --------------- Transmit Ports - TX Driver and OOB signalling --------------
        TXN0_OUT                        =>      TILE1_TXN0_OUT,
        TXN1_OUT                        =>      TILE1_TXN1_OUT,
        TXP0_OUT                        =>      TILE1_TXP0_OUT,
        TXP1_OUT                        =>      TILE1_TXP1_OUT,
        -------- Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
        TXENPMAPHASEALIGN0_IN           =>      TILE1_TXENPMAPHASEALIGN0_IN,
        TXENPMAPHASEALIGN1_IN           =>      TILE1_TXENPMAPHASEALIGN1_IN,
        TXPMASETPHASE0_IN               =>      TILE1_TXPMASETPHASE0_IN,
        TXPMASETPHASE1_IN               =>      TILE1_TXPMASETPHASE1_IN,
        -------------------- Transmit Ports - polarity  ----------------------------
        TXPOLARITY0                     =>      TILE1_TXPOLARITY0,
        TXPOLARITY1                     =>      TILE1_TXPOLARITY1,
        ----------------- Transmit Ports - TX Ports for PCI Express ----------------
        TXELECIDLE0_IN                  =>      TILE1_TXELECIDLE0_IN,
        TXELECIDLE1_IN                  =>      TILE1_TXELECIDLE1_IN
    );
end generate;  

GEN_SWAP1: if (CH23_SWAP) generate
    --_________________________________________________________________________
    --_________________________________________________________________________
    --TILE1  (Location)

    tile1_rocketio_wrapper_i : ROCKETIO_WRAPPER_TILE
    generic map
    (
        -- Simulation attributes
        TILE_SIM_MODE                => WRAPPER_SIM_MODE,
        TILE_SIM_GTXRESET_SPEEDUP    => WRAPPER_SIM_GTXRESET_SPEEDUP,
        TILE_SIM_PLL_PERDIV2         => WRAPPER_SIM_PLL_PERDIV2,

        -- Channel bonding attributes
        TILE_CHAN_BOND_MODE_0        => "SLAVE",
        TILE_CHAN_BOND_LEVEL_0       => 1,

        TILE_CHAN_BOND_MODE_1        => "MASTER",
        TILE_CHAN_BOND_LEVEL_1       => 2
    )
    port map
    (
        ------------------------ Loopback and Powerdown Ports ----------------------
        LOOPBACK0_IN                    =>      TILE1_LOOPBACK1_IN,
        LOOPBACK1_IN                    =>      TILE1_LOOPBACK0_IN,
        RXPOWERDOWN0_IN                 =>      TILE1_RXPOWERDOWN1_IN,
        RXPOWERDOWN1_IN                 =>      TILE1_RXPOWERDOWN0_IN,
        TXPOWERDOWN0_IN                 =>      TILE1_TXPOWERDOWN1_IN,
        TXPOWERDOWN1_IN                 =>      TILE1_TXPOWERDOWN0_IN,
        ----------------------- Receive Ports - 8b10b Decoder ----------------------
        RXCHARISCOMMA0_OUT              =>      tile1_rxchariscomma1_i,
        RXCHARISCOMMA1_OUT              =>      tile1_rxchariscomma0_i,
        RXCHARISK0_OUT                  =>      tile1_rxcharisk1_i,
        RXCHARISK1_OUT                  =>      tile1_rxcharisk0_i,
        RXDISPERR0_OUT                  =>      tile1_rxdisperr1_i,
        RXDISPERR1_OUT                  =>      tile1_rxdisperr0_i,
        RXNOTINTABLE0_OUT               =>      tile1_rxnotintable1_i,
        RXNOTINTABLE1_OUT               =>      tile1_rxnotintable0_i,
        RXRUNDISP0_OUT                  =>      tile1_rxrundisp1_i,
        RXRUNDISP1_OUT                  =>      tile1_rxrundisp0_i,
        ------------------- Receive Ports - Channel Bonding Ports ------------------
        RXCHANBONDSEQ0_OUT              =>      tile1_rxchanbondseq1_i,
        RXCHANBONDSEQ1_OUT              =>      tile1_rxchanbondseq0_i,
        RXCHBONDI0_IN                   =>      tile1_rxchbondo0_i,
        RXCHBONDI1_IN                   =>      tied_to_ground_vec_i(3 downto 0),
        RXCHBONDO0_OUT                  =>      tile1_rxchbondo1_i,
        RXCHBONDO1_OUT                  =>      tile1_rxchbondo0_i,
        RXENCHANSYNC0_IN                =>      TILE1_RXENCHANSYNC1_IN,
        RXENCHANSYNC1_IN                =>      TILE1_RXENCHANSYNC0_IN,
        ------------------- Receive Ports - Clock Correction Ports -----------------
        RXCLKCORCNT0_OUT                =>      tile1_rxclkcorcnt1_i,
        RXCLKCORCNT1_OUT                =>      tile1_rxclkcorcnt0_i,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        RXBYTEISALIGNED0_OUT            =>      TILE1_RXBYTEISALIGNED1_OUT,
        RXBYTEISALIGNED1_OUT            =>      TILE1_RXBYTEISALIGNED0_OUT,
        RXBYTEREALIGN0_OUT              =>      TILE1_RXBYTEREALIGN1_OUT,
        RXBYTEREALIGN1_OUT              =>      TILE1_RXBYTEREALIGN0_OUT,
        RXCOMMADET0_OUT                 =>      TILE1_RXCOMMADET1_OUT,
        RXCOMMADET1_OUT                 =>      TILE1_RXCOMMADET0_OUT,
        RXENMCOMMAALIGN0_IN             =>      TILE1_RXENMCOMMAALIGN1_IN,
        RXENMCOMMAALIGN1_IN             =>      TILE1_RXENMCOMMAALIGN0_IN,
        RXENPCOMMAALIGN0_IN             =>      TILE1_RXENPCOMMAALIGN1_IN,
        RXENPCOMMAALIGN1_IN             =>      TILE1_RXENPCOMMAALIGN0_IN,
        ------------------- Receive Ports - RX Data Path interface -----------------
        RXDATA0_OUT                     =>      tile1_rxdata1_i,
        RXDATA1_OUT                     =>      tile1_rxdata0_i,
        RXRECCLK0_OUT                   =>      tile1_rxrecclk1_i,
        RXRECCLK1_OUT                   =>      tile1_rxrecclk0_i,
        RXRESET0_IN                     =>      tile1_rxreset1_i,
        RXRESET1_IN                     =>      tile1_rxreset0_i,
        RXUSRCLK0_IN                    =>      tile1_rxrecclk0_bufg_i,
        RXUSRCLK1_IN                    =>      tile1_rxrecclk0_bufg_i,
        RXUSRCLK20_IN                   =>      tile1_rxrecclk0_bufg_i,
        RXUSRCLK21_IN                   =>      tile1_rxrecclk0_bufg_i,
        ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        RXCDRRESET0_IN                  =>      TILE1_RXCDRRESET1_IN,
        RXCDRRESET1_IN                  =>      TILE1_RXCDRRESET0_IN,
        RXELECIDLE0_OUT                 =>      TILE1_RXELECIDLE1_OUT,
        RXELECIDLE1_OUT                 =>      TILE1_RXELECIDLE0_OUT,
        RXN0_IN                         =>      TILE1_RXN1_IN,
        RXN1_IN                         =>      TILE1_RXN0_IN,
        RXP0_IN                         =>      TILE1_RXP1_IN,
        RXP1_IN                         =>      TILE1_RXP0_IN,
        -------- Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
        RXBUFRESET0_IN                  =>      tile1_rxbufreset1_i,
        RXBUFRESET1_IN                  =>      tile1_rxbufreset0_i,
        RXBUFSTATUS0_OUT                =>      tile1_rxbufstatus1_i,
        RXBUFSTATUS1_OUT                =>      tile1_rxbufstatus0_i,
        RXCHANISALIGNED0_OUT            =>      tile1_rxchanisaligned1_i,
        RXCHANISALIGNED1_OUT            =>      tile1_rxchanisaligned0_i,
        RXCHANREALIGN0_OUT              =>      tile1_rxchanrealign1_i,
        RXCHANREALIGN1_OUT              =>      tile1_rxchanrealign0_i,
        --------------- Receive Ports - RX Loss-of-sync State Machine --------------
        RXLOSSOFSYNC0_OUT               =>      tile1_rxlossofsync1_i,
        RXLOSSOFSYNC1_OUT               =>      tile1_rxlossofsync0_i,
        -------------- Receive Ports - polarity  -----------------------------------
        RXPOLARITY0                     =>      TILE1_RXPOLARITY1,
        RXPOLARITY1                     =>      TILE1_RXPOLARITY0,
        -------------- Receive Ports - RX Pipe Control for PCI Express -------------
        RXVALID0_OUT                    =>      tile1_rxvalid1_i,
        RXVALID1_OUT                    =>      tile1_rxvalid0_i,
        ------------- Shared Ports - Dynamic Reconfiguration Port (DRP) ------------
        DADDR_IN                        =>      TILE1_DADDR_IN,
        DCLK_IN                         =>      TILE1_DCLK_IN,
        DEN_IN                          =>      TILE1_DEN_IN,
        DI_IN                           =>      TILE1_DI_IN,
        DO_OUT                          =>      TILE1_DO_OUT,
        DRDY_OUT                        =>      TILE1_DRDY_OUT,
        DWE_IN                          =>      TILE1_DWE_IN,
        --------------------- Shared Ports - Tile and PLL Ports --------------------
        CLKIN_IN                        =>      TILE1_CLKIN_IN,
        GTXRESET_IN                     =>      TILE1_GTXRESET_IN,
        PLLLKDET_OUT                    =>      TILE1_PLLLKDET_OUT,
        REFCLKOUT_OUT                   =>      TILE1_REFCLKOUT_OUT,
        RESETDONE0_OUT                  =>      tile1_resetdone1_i,
        RESETDONE1_OUT                  =>      tile1_resetdone0_i,
        ---------------- Transmit Ports - 8b10b Encoder Control Ports --------------
        TXCHARISK0_IN                   =>      TILE1_TXCHARISK1_IN,
        TXCHARISK1_IN                   =>      TILE1_TXCHARISK0_IN,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        TXDATA0_IN                      =>      TILE1_TXDATA1_IN,
        TXDATA1_IN                      =>      TILE1_TXDATA0_IN,
        TXRESET0_IN                     =>      TILE1_TXRESET1_IN,
        TXRESET1_IN                     =>      TILE1_TXRESET0_IN,
        TXUSRCLK0_IN                    =>      TILE1_TXUSRCLK1_IN,
        TXUSRCLK1_IN                    =>      TILE1_TXUSRCLK0_IN,
        TXUSRCLK20_IN                   =>      TILE1_TXUSRCLK21_IN,
        TXUSRCLK21_IN                   =>      TILE1_TXUSRCLK20_IN,
        --------------- Transmit Ports - TX Driver and OOB signalling --------------
        TXN0_OUT                        =>      TILE1_TXN1_OUT,
        TXN1_OUT                        =>      TILE1_TXN0_OUT,
        TXP0_OUT                        =>      TILE1_TXP1_OUT,
        TXP1_OUT                        =>      TILE1_TXP0_OUT,
        -------- Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
        TXENPMAPHASEALIGN0_IN           =>      TILE1_TXENPMAPHASEALIGN1_IN,
        TXENPMAPHASEALIGN1_IN           =>      TILE1_TXENPMAPHASEALIGN0_IN,
        TXPMASETPHASE0_IN               =>      TILE1_TXPMASETPHASE1_IN,
        TXPMASETPHASE1_IN               =>      TILE1_TXPMASETPHASE0_IN,
        -------------------- Transmit Ports - polarity  ----------------------------
        TXPOLARITY0                     =>      TILE1_TXPOLARITY1,
        TXPOLARITY1                     =>      TILE1_TXPOLARITY0,
        ----------------- Transmit Ports - TX Ports for PCI Express ----------------
        TXELECIDLE0_IN                  =>      TILE1_TXELECIDLE1_IN,
        TXELECIDLE1_IN                  =>      TILE1_TXELECIDLE0_IN
    );
end generate;  

    --_________________________________________________________________________
    --_________________________________________________________________________
    tile1_rxrecclk0_bufg0_i : BUFG
    port map
    (
        I                               =>      tile1_rxrecclk0_i,
        O                               =>      tile1_rxrecclk0_bufg_i
    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --TILE1 GTP0
    tile1_gtp0_cc_2b_1skp_i : CC_2B_1SKP
    generic map
    (
        CC_CHAR                      => x"1c",
        ALIGN_CHAR                   => x"7c",
        CHAN_BOND_MODE               => "MASTER",
        ALIGN_PARALLEL_CHECK         => '1'
    )
    port map
    (
        -- Write Interface on the RXRECCLK
        GT_RXDATA                       =>      tile1_rxdata0_i,
        GT_RXCHARISK                    =>      tile1_rxcharisk0_i,
        GT_RXCHARISCOMMA                =>      tile1_rxchariscomma0_i,
        GT_RXRUNDISP                    =>      tile1_rxrundisp0_i,
        GT_RXNOTINTABLE                 =>      tile1_rxnotintable0_i,
        GT_RXDISPERR                    =>      tile1_rxdisperr0_i,
        GT_RXBUFSTATUS                  =>      tile1_rxbufstatus0_i,
        GT_RXCLKCORCNT                  =>      tile1_rxclkcorcnt0_i,
        GT_RXCHANBONDSEQ                =>      tile1_rxchanbondseq0_i,
        GT_RXCHANISALIGNED              =>      tile1_rxchanisaligned0_i,
        GT_RXCHANREALIGN                =>      tile1_rxchanrealign0_i,
        GT_RXLOSSOFSYNC                 =>      tile1_rxlossofsync0_i,
        GT_RXVALID                      =>      tile1_rxvalid0_i,
        GT_RXUSRCLK2                    =>      tile1_rxrecclk0_bufg_i,

        -- Read Interface on the RXUSRCLK2
        USER_RXDATA                     =>      TILE1_RXDATA0_OUT,
        USER_RXCHARISK                  =>      TILE1_RXCHARISK0_OUT,
        USER_RXCHARISCOMMA              =>      TILE1_RXCHARISCOMMA0_OUT,
        USER_RXRUNDISP                  =>      open,
        USER_RXNOTINTABLE               =>      TILE1_RXNOTINTABLE0_OUT,
        USER_RXDISPERR                  =>      TILE1_RXDISPERR0_OUT,
        USER_RXBUFSTATUS                =>      TILE1_RXBUFSTATUS0_OUT,
        USER_RXCLKCORCNT                =>      TILE1_RXCLKCORCNT0_OUT,
        USER_RXCHANBONDSEQ              =>      TILE1_RXCHANBONDSEQ0_OUT,
        USER_RXCHANISALIGNED            =>      TILE1_RXCHANISALIGNED0_OUT,
        USER_RXCHANREALIGN              =>      TILE1_RXCHANREALIGN0_OUT,
        USER_RXLOSSOFSYNC               =>      TILE1_RXLOSSOFSYNC0_OUT,
        USER_RXVALID                    =>      open,
        USER_RXUSRCLK2                  =>      TILE1_RXUSRCLK20_IN,

        -- Status and reset signals
        RESET                           =>      tile1_gtp0_cc_2b_1skp_reset_i,
        CCI                             =>      tied_to_ground_vec_i(6 downto 0),
        CCO                             =>      tile1_gtp0_cc_2b_1skp_cco_i
    );


    -- Reset logic
    tile1_gtp0_cc_2b_1skp_reset_i <= (not(tile0_resetdone0_i
                                           and tile0_resetdone1_i
                                           and tile1_resetdone0_i
                                           and tile1_resetdone1_i))
                                            or tile1_rxreset0_i or tile1_rxbufreset0_i;

    TILE1_RESETDONE0_OUT <= tile1_resetdone0_i;
    tile1_rxreset0_i <= TILE1_RXRESET0_IN;
    tile1_rxbufreset0_i <= TILE1_RXBUFRESET0_IN;


    --_________________________________________________________________________
    --_________________________________________________________________________
    --TILE1 GTP1
    tile1_gtp1_cc_2b_1skp_i : CC_2B_1SKP
    generic map
    (
        CC_CHAR                      => x"1c",
        ALIGN_CHAR                   => x"7c",
        CHAN_BOND_MODE               => "SLAVE",
        ALIGN_PARALLEL_CHECK         => '1'
    )
    port map
    (
        -- Write Interface on the RXRECCLK
        GT_RXDATA                       =>      tile1_rxdata1_i,
        GT_RXCHARISK                    =>      tile1_rxcharisk1_i,
        GT_RXCHARISCOMMA                =>      tile1_rxchariscomma1_i,
        GT_RXRUNDISP                    =>      tile1_rxrundisp1_i,
        GT_RXNOTINTABLE                 =>      tile1_rxnotintable1_i,
        GT_RXDISPERR                    =>      tile1_rxdisperr1_i,
        GT_RXBUFSTATUS                  =>      tile1_rxbufstatus1_i,
        GT_RXCLKCORCNT                  =>      tile1_rxclkcorcnt1_i,
        GT_RXCHANBONDSEQ                =>      tile1_rxchanbondseq1_i,
        GT_RXCHANISALIGNED              =>      tile1_rxchanisaligned1_i,
        GT_RXCHANREALIGN                =>      tile1_rxchanrealign1_i,
        GT_RXLOSSOFSYNC                 =>      tile1_rxlossofsync1_i,
        GT_RXVALID                      =>      tile1_rxvalid1_i,
        GT_RXUSRCLK2                    =>      tile1_rxrecclk0_bufg_i,

        -- Read Interface on the RXUSRCLK2
        USER_RXDATA                     =>      TILE1_RXDATA1_OUT,
        USER_RXCHARISK                  =>      TILE1_RXCHARISK1_OUT,
        USER_RXCHARISCOMMA              =>      TILE1_RXCHARISCOMMA1_OUT,
        USER_RXRUNDISP                  =>      open,
        USER_RXNOTINTABLE               =>      TILE1_RXNOTINTABLE1_OUT,
        USER_RXDISPERR                  =>      TILE1_RXDISPERR1_OUT,
        USER_RXBUFSTATUS                =>      TILE1_RXBUFSTATUS1_OUT,
        USER_RXCLKCORCNT                =>      TILE1_RXCLKCORCNT1_OUT,
        USER_RXCHANBONDSEQ              =>      TILE1_RXCHANBONDSEQ1_OUT,
        USER_RXCHANISALIGNED            =>      TILE1_RXCHANISALIGNED1_OUT,
        USER_RXCHANREALIGN              =>      TILE1_RXCHANREALIGN1_OUT,
        USER_RXLOSSOFSYNC               =>      TILE1_RXLOSSOFSYNC1_OUT,
        USER_RXVALID                    =>      open,
        USER_RXUSRCLK2                  =>      TILE1_RXUSRCLK21_IN,

        -- Status and reset signals
        RESET                           =>      tied_to_ground_i,
        CCI                             =>      tile1_gtp0_cc_2b_1skp_cco_i,
        CCO                             =>      open
    );

    TILE1_RESETDONE1_OUT <= tile1_resetdone1_i;
    tile1_rxreset1_i <= TILE1_RXRESET1_IN;
    tile1_rxbufreset1_i <= TILE1_RXBUFRESET1_IN;

end RTL;
