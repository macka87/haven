/*
 * IB_TRANSFORMER_8_64.sv: IB_TRANSFORMER System Verilog envelope
 * Copyright (C) 2008 CESNET
 * Author(s): Tomas Malek <tomalek@liberouter.org>
 *
 * Redistribution and use in source and binary forms, with or without
 * modification, are permitted provided that the following conditions
 * are met:
 * 1. Redistributions of source code must retain the above copyright
 *    notice, this list of conditions and the following disclaimer.
 * 2. Redistributions in binary form must reproduce the above copyright
 *    notice, this list of conditions and the following disclaimer in
 *    the documentation and/or other materials provided with the
 *    distribution.
 * 3. Neither the name of the Company nor the names of its contributors
 *    may be used to endorse or promote products derived from this
 *    software without specific prior written permission.
 *
 * This software is provided ``as is'', and any express or implied
 * warranties, including, but not limited to, the implied warranties of
 * merchantability and fitness for a particular purpose are disclaimed.
 * In no event shall the company or contributors be liable for any
 * direct, indirect, incidental, special, exemplary, or consequential
 * damages (including, but not limited to, procurement of substitute
 * goods or services; loss of use, data, or profits; or business
 * interruption) however caused and on any theory of liability, whether
 * in contract, strict liability, or tort (including negligence or
 * otherwise) arising in any way out of the use of this software, even
 * if advised of the possibility of such damage.
 *
 * $Id: ib_transformer_8_64.sv 1899 2008-03-26 15:52:13Z tomalek $
 *
 * TODO:
 *
 */
 
module IB_TRANSFORMER_8_64_SV (
   input logic CLK,
   input logic RESET,
   iIB64.rx UP_IN,
   iIB64.tx UP_OUT,
   iIB8.tx DOWN_OUT,
   iIB8.rx DOWN_IN);

   IB_TRANSFORMER TRANSFORMER_INST (
      // Common Interface
      .CLK               (CLK),
      .RESET             (RESET),

      // UP port
      .UP_IN_DATA         (UP_IN.DATA),         
      .UP_IN_SOF_N        (UP_IN.SOF_N),        
      .UP_IN_EOF_N        (UP_IN.EOF_N),        
      .UP_IN_SRC_RDY_N    (UP_IN.SRC_RDY_N),    
      .UP_IN_DST_RDY_N    (UP_IN.DST_RDY_N),    
                                              
      .UP_OUT_DATA        (UP_OUT.DATA),        
      .UP_OUT_SOF_N       (UP_OUT.SOF_N),       
      .UP_OUT_EOF_N       (UP_OUT.EOF_N),       
      .UP_OUT_SRC_RDY_N   (UP_OUT.SRC_RDY_N),   
      .UP_OUT_DST_RDY_N   (UP_OUT.DST_RDY_N),   
                                              
      // DOWN port        
      .DOWN_OUT_DATA      (DOWN_OUT.DATA),      
      .DOWN_OUT_SOF_N     (DOWN_OUT.SOF_N),     
      .DOWN_OUT_EOF_N     (DOWN_OUT.EOF_N),     
      .DOWN_OUT_SRC_RDY_N (DOWN_OUT.SRC_RDY_N), 
      .DOWN_OUT_DST_RDY_N (DOWN_OUT.DST_RDY_N), 
                                              
      .DOWN_IN_DATA       (DOWN_IN.DATA),       
      .DOWN_IN_SOF_N      (DOWN_IN.SOF_N),      
      .DOWN_IN_EOF_N      (DOWN_IN.EOF_N),      
      .DOWN_IN_SRC_RDY_N  (DOWN_IN.SRC_RDY_N),  
      .DOWN_IN_DST_RDY_N  (DOWN_IN.DST_RDY_N)        
);

endmodule : IB_TRANSFORMER_8_64_SV



