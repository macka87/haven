/* *****************************************************************************
 * Project Name: HAVEN
 * File Name:    sv_alu_seq_pkg.sv
 * Description:  OVM ALU Sequence Package
 * Authors:      Michaela Belesova <xbeles00@stud.fit.vutbr.cz>,
 *               Marcela Simkova <isimkova@fit.vutbr.cz> 
 * Date:         26.9.2012
 * ************************************************************************** */

package sv_alu_seq_pkg;

endpackage