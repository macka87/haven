--
-- input.vhd : Internal Bus Switch Input entity
-- Copyright (C) 2008 CESNET
-- Author(s): Tomas Malek <tomalek@liberouter.org>
--
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above copyright
--    notice, this list of conditions and the following disclaimer in
--    the documentation and/or other materials provided with the
--    distribution.
-- 3. Neither the name of the Company nor the names of its contributors
--    may be used to endorse or promote products derived from this
--    software without specific prior written permission.
--
-- This software is provided ``as is'', and any express or implied
-- warranties, including, but not limited to, the implied warranties of
-- merchantability and fitness for a particular purpose are disclaimed.
-- In no event shall the company or contributors be liable for any
-- direct, indirect, incidental, special, exemplary, or consequential
-- damages (including, but not limited to, procurement of substitute
-- goods or services; loss of use, data, or profits; or business
-- interruption) however caused and on any theory of liability, whether
-- in contract, strict liability, or tort (including negligence or
-- otherwise) arising in any way out of the use of this software, even
-- if advised of the possibility of such damage.
--
-- $Id$
--
-- TODO:
-- 

library IEEE;
use IEEE.std_logic_1164.all;

-- ----------------------------------------------------------------------------
--                    ENTITY DECLARATION -- IB Switch Input                  --
-- ----------------------------------------------------------------------------
      
entity IB_SWITCH_INPUT is 
   generic(
      -- Data Width (1-128)
      DATA_WIDTH   : integer:= 64;
      -- Port 1 Address Space
      PORT1_BASE   : std_logic_vector(31 downto 0) := X"11111111";
      PORT1_LIMIT  : std_logic_vector(31 downto 0) := X"11111111";
      -- Port 2 Address Space
      PORT2_BASE   : std_logic_vector(31 downto 0) := X"22222222"; 
      PORT2_LIMIT  : std_logic_vector(31 downto 0) := X"22222222"   
   ); 
   port (
      -- Common interface -----------------------------------------------------
      CLK            : in std_logic;  
      RESET          : in std_logic;  

      -- Upstream Port #0 -----------------------------------------------------
      -- input ifc --            
      IN0_DATA      : in  std_logic_vector(DATA_WIDTH-1 downto 0);
      IN0_SOF_N     : in  std_logic;
      IN0_EOF_N     : in  std_logic;
      IN0_SRC_RDY_N : in  std_logic;
      IN0_DST_RDY_N : out std_logic;

      -- output ifc --
      OUT0_DATA      : out std_logic_vector(DATA_WIDTH-1 downto 0);
      OUT0_SOF_N     : out std_logic;
      OUT0_EOF_N     : out std_logic;
      OUT0_WR        : out std_logic;
      OUT0_FULL      : in  std_logic;      

      OUT0_REQ_VEC   : out std_logic_vector(2 downto 0);
      OUT0_REQ_WE    : out std_logic;      

      -- Downstream Port #1 ---------------------------------------------------
      -- input ifc --            
      IN1_DATA      : in  std_logic_vector(DATA_WIDTH-1 downto 0);
      IN1_SOF_N     : in  std_logic;
      IN1_EOF_N     : in  std_logic;
      IN1_SRC_RDY_N : in  std_logic;
      IN1_DST_RDY_N : out std_logic;
        
      -- output ifc --
      OUT1_DATA      : out std_logic_vector(DATA_WIDTH-1 downto 0);
      OUT1_SOF_N     : out std_logic;
      OUT1_EOF_N     : out std_logic;
      OUT1_WR        : out std_logic;
      OUT1_FULL      : in  std_logic;    

      OUT1_REQ_VEC   : out std_logic_vector(2 downto 0);
      OUT1_REQ_WE    : out std_logic;      
      
      -- Downstream Port #2 ---------------------------------------------------
      -- input ifc --            
      IN2_DATA      : in  std_logic_vector(DATA_WIDTH-1 downto 0);
      IN2_SOF_N     : in  std_logic;
      IN2_EOF_N     : in  std_logic;
      IN2_SRC_RDY_N : in  std_logic;
      IN2_DST_RDY_N : out std_logic;

      -- output ifc --
      OUT2_DATA      : out std_logic_vector(DATA_WIDTH-1 downto 0);
      OUT2_SOF_N     : out std_logic;
      OUT2_EOF_N     : out std_logic;
      OUT2_WR        : out std_logic;
      OUT2_FULL      : in  std_logic;          
      
      OUT2_REQ_VEC   : out std_logic_vector(2 downto 0);
      OUT2_REQ_WE    : out std_logic          
   );
end IB_SWITCH_INPUT;



