/* *****************************************************************************
 * Project Name: NetCOPE Adder Functional Verification
 * File Name:    test_pkg.sv - test package
 * Description:  Definition of constants and parameters 
 * Author:       Marcela Simkova <xsimko03@stud.fit.vutbr.cz> 
 * Date:         27.2.2011 
 * ************************************************************************** */ 

package test_pkg;
   
   import math_pkg::*;       
   
   // VERIFICATION FRAMEWORK
   int FRAMEWORK  = 0;                         // 0 = software framework
                                               // 1 = sw/hw framework      
   // DUT GENERICS
   parameter DATA_WIDTH = 128;                 // FrameLink data width
   parameter DREM_WIDTH = log2(DATA_WIDTH/8);  // drem width
   
   // CLOCKS AND RESETS
   parameter CLK_PERIOD = 10ns;
   parameter RESET_TIME = 10*CLK_PERIOD;

   // TRANSACTION FORMAT 
   int GENERATOR_FL_FRAME_COUNT     = 1;       // frame parts
   int GENERATOR_FL_PART_SIZE_MAX[] = '{36};   // maximal size of part
   int GENERATOR_FL_PART_SIZE_MIN[] = '{1};    // minimal size of part     
   
   // SOFTWARE DRIVER PARAMETERS 
   // Enable/Disable weights of "delay between transactions" 
   parameter DRIVER_BT_DELAY_EN_WT  = 0;       
   parameter DRIVER_BT_DELAY_DI_WT  = 5;
   // Low/High limit of "delay between transactions" value
   parameter DRIVER_BT_DELAY_LOW    = 0;
   parameter DRIVER_BT_DELAY_HIGH   = 10;
   // Enable/Disable weights of "delays inside transaction"
   parameter DRIVER_IT_DELAY_EN_WT  = 0;
   parameter DRIVER_IT_DELAY_DI_WT  = 5;
   // Low/High limit of "delay inside transaction" values
   parameter DRIVER_IT_DELAY_LOW    = 0;
   parameter DRIVER_IT_DELAY_HIGH   = 10;

   // TEST PARAMETERS
   parameter TRANSACTION_COUT = 1;            // Count of transactions

endpackage
