/* *****************************************************************************
 * Project Name: HAVEN - Genetic Algorithm
 * File Name:    sv_alu_seq_pkg.sv
 * Description:  UVM ALU Sequence Package
 * Authors:      Marcela Simkova <isimkova@fit.vutbr.cz> 
 * Date:         19.4.2013
 * ************************************************************************** */

 package sv_alu_seq_pkg;

   // Standard UVM import & include
   import uvm_pkg::*;
   `include "uvm_macros.svh"
  
   // Package imports
   import sv_alu_param_pkg::*;
   //import sv_basic_ga_pkg::*;
  
   // Includes  !! svh !!
   /*`include "alu_chromosome.sv"
   `include "haven_sequence_item.sv"
   `include "haven_input_transaction.sv"
   `include "haven_output_transaction.sv"
   `include "alu_input_transaction.sv"
   `include "alu_output_transaction.sv"
   `include "alu_sequence.sv"
   `include "alu_sequencer.sv" */
  
 endpackage