/*
 * fl_fifo_ifc.sv: FrameLink FIFO Control Interface
 * Copyright (C) 2008 CESNET
 * Author(s): Marek Santa <xsanta06@stud.fit.vutbr.cz>
 *
 * Redistribution and use in source and binary forms, with or without
 * modification, are permitted provided that the following conditions
 * are met:
 * 1. Redistributions of source code must retain the above copyright
 *    notice, this list of conditions and the following disclaimer.
 * 2. Redistributions in binary form must reproduce the above copyright
 *    notice, this list of conditions and the following disclaimer in
 *    the documentation and/or other materials provided with the
 *    distribution.
 * 3. Neither the name of the Company nor the names of its contributors
 *    may be used to endorse or promote products derived from this
 *    software without specific prior written permission.
 *
 * This software is provided ``as is'', and any express or implied
 * warranties, including, but not limited to, the implied warranties of
 * merchantability and fitness for a particular purpose are disclaimed.
 * In no event shall the company or contributors be liable for any
 * direct, indirect, incidental, special, exemplary, or consequential
 * damages (including, but not limited to, procurement of substitute
 * goods or services; loss of use, data, or profits; or business
 * interruption) however caused and on any theory of liability, whether
 * in contract, strict liability, or tort (including negligence or
 * otherwise) arising in any way out of the use of this software, even
 * if advised of the possibility of such damage.
 *
 * $Id: fl_fifo_ifc.sv 5883 2008-10-10 22:39:52Z xsanta06 $
 *
 * TODO:
 *
 */
 

// ----------------------------------------------------------------------------
//                 FrameLink FIFO Control Interface declaration
// ----------------------------------------------------------------------------

// -- FrameLink FIFO Control Interface ----------------------------------------
interface iFrameLinkFifo #(STATUS_WIDTH = 8) (input logic CLK, RESET);  
  // Control Interface
  logic LSTBLK                    ;   // Last block detection
  logic [STATUS_WIDTH-1:0] STATUS ;   // MSBs of exact number of free items in the FIFO
  logic EMPTY                     ;   // FIFO is empty
  logic FULL                      ;   // FIFO is full
  logic FRAME_RDY                 ;   // At least one whole frame is in the FIFO
    

  // Clocking blocks  
  clocking ctrl_cb @(posedge CLK);
    input  LSTBLK, STATUS, EMPTY, FULL, FRAME_RDY;
  endclocking: ctrl_cb;

  // Control Modport
  modport ctrl (output  LSTBLK,
                output  STATUS,
                output  EMPTY,
                output  FULL,
                output  FRAME_RDY
               );
  
  modport ctrl_tb (clocking ctrl_cb);

endinterface : iFrameLinkFifo
