-- fl_watch_lb.vhd: Frame Link watch local bus cover.
-- Copyright (C) 2006 CESNET
-- Author(s): Viktor Pus <pus@liberouter.org>
--            Lukas Solanka <solanka@liberouter.org>
--
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above copyright
--    notice, this list of conditions and the following disclaimer in
--    the documentation and/or other materials provided with the
--    distribution.
-- 3. Neither the name of the Company nor the names of its contributors
--    may be used to endorse or promote products derived from this
--    software without specific prior written permission.
--
-- This software is provided ``as is'', and any express or implied
-- warranties, including, but not limited to, the implied warranties of
-- merchantability and fitness for a particular purpose are disclaimed.
-- In no event shall the company or contributors be liable for any
-- direct, indirect, incidental, special, exemplary, or consequential
-- damages (including, but not limited to, procurement of substitute
-- goods or services; loss of use, data, or profits; or business
-- interruption) however caused and on any theory of liability, whether
-- in contract, strict liability, or tort (including negligence or
-- otherwise) arising in any way out of the use of this software, even
-- if advised of the possibility of such damage.
--
-- $Id$
--

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

-- Library with MI32 interface definition
use work.lb_pkg.all;

-- library containing log2 function
use work.math_pack.all;

-- ----------------------------------------------------------------------------
--                            Entity declaration
-- ----------------------------------------------------------------------------
entity FL_WATCH_LB is
   generic(
      INTERFACES     : integer := 1;  -- At least 1
      CNTR_WIDTH     : integer := 32;
      PIPELINE_LEN   : integer := 1;   -- At least 1
      GUARD          : boolean := true;
      HEADER         : boolean := true;
      FOOTER         : boolean := true;

      -- Local bus
      BASE_ADDR      : integer;   -- base address 
      ADDR_WIDTH     : integer;   -- address width
      FREQUENCY      : integer := 100 -- frequency
   );
   port(
      CLK            : in  std_logic;
      RESET          : in  std_logic;

      SOF_N          : in std_logic_vector(INTERFACES-1 downto 0);
      EOF_N          : in std_logic_vector(INTERFACES-1 downto 0);
      SOP_N          : in std_logic_vector(INTERFACES-1 downto 0);
      EOP_N          : in std_logic_vector(INTERFACES-1 downto 0);
      DST_RDY_N      : in std_logic_vector(INTERFACES-1 downto 0);
      SRC_RDY_N      : in std_logic_vector(INTERFACES-1 downto 0);

      -- Local bus signals
      LBCLK       : in    std_logic; 
      LBFRAME     : in    std_logic; -- Frame
      LBHOLDA     : out   std_logic; -- Hold Ack (HOLDA), active LOW
      LBAD        : inout std_logic_vector(15 downto 0); -- Address/Data
      LBAS        : in    std_logic; -- Adress strobe
      LBRW        : in    std_logic;
      LBRDY       : out   std_logic; -- Ready, active LOW
      LBLAST      : in    std_logic
   );
end entity FL_WATCH_LB;


-- ----------------------------------------------------------------------------
--                               Architecture
-- ----------------------------------------------------------------------------
architecture full of FL_WATCH_LB is
   -- MI32 connection
   signal mi : t_mi32;
begin

   FL_WATCH_MI_U: entity work.FL_WATCH
      generic map (
         INTERFACES     => INTERFACES,
         CNTR_WIDTH     => CNTR_WIDTH,
         PIPELINE_LEN   => PIPELINE_LEN,
         GUARD          => GUARD,
         HEADER         => HEADER,
         FOOTER         => FOOTER
      )
      port map (
         CLK            => CLK,
         RESET          => RESET,
   
         SOF_N          => SOF_N,
         EOF_N          => EOF_N,
         SOP_N          => SOP_N,
         EOP_N          => EOP_N,
         DST_RDY_N      => DST_RDY_N,
         SRC_RDY_N      => SRC_RDY_N,
   
         MI             => mi
      );
   
   mi.addr(31 downto ADDR_WIDTH) <= (others => '0');
   mi.be <= (others => '1');
   
   LB_CONNECT_U: entity work.lb_connect
      generic map (
         BASE_ADDR  => BASE_ADDR,
         ADDR_WIDTH => ADDR_WIDTH,
         FREQUENCY  => FREQUENCY
      )
      port map (
         -- Control signals
         RESET             => RESET,
   
         -- LB signals
         LBCLK       => LBCLK,
         LBFRAME     => LBFRAME,
         LBHOLDA     => LBHOLDA,
         LBAD        => LBAD,
         LBAS        => LBAS,
         LBRW        => LBRW,
         LBRDY       => LBRDY,
         LBLAST      => LBLAST,
   
         -- Address decoder interface
         CLK         => CLK,
         ADC_RD      => mi.rd,
         ADC_WR      => mi.wr,
         ADC_ADDR    => mi.addr(ADDR_WIDTH - 1 downto 0),
         ADC_DI      => mi.dwr,
         ADC_DO      => mi.drd,
         ADC_DRDY    => mi.drdy
      );

end architecture full;


