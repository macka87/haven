/* *****************************************************************************
 * Project Name: HAVEN
 * File Name:    alu_general_settings.sv
 * Description:  Changeable settings
 * Authors:      Michaela Belesova <xbeles00@stud.fit.vutbr.cz>,
 *               Marcela Simkova <isimkova@fit.vutbr.cz> 
 * Date:         13.9.2012
 * ************************************************************************** */
 
 package alu_general_settings_pkg;
 
   // DUT GENERICS
   parameter DATA_WIDTH     = 8;
   
   // CLOCK
   parameter CLK_PERIOD     = 10ns;
   
 endpackage