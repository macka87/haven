/* *****************************************************************************
 * Project Name: Software Framework for Functional Verification
 * File Name:    sv_basic_comp_pkg.sv
 * Description:  SystemVerilog Basic Verification Components 
 * Author:       Marcela Simkova <xsimko03@stud.fit.vutbr.cz> 
 * Date:         27.2.2011 
 * ************************************************************************** */

package sv_basic_comp_pkg; 
   import sv_types_pkg::*; // Import package of user defined types 

  `include "transaction.sv"
  `include "netcope_transaction.sv"
  `include "generator.sv"
  `include "input_cbs.sv"
  `include "input_controller.sv"
  `include "gen_input_controller.sv"    
  `include "driver.sv"
  `include "sender.sv"
  `include "dpi/input_wrapper.sv"
  `include "dpi/output_wrapper.sv"
  `include "sorter.sv"
  `include "output_cbs.sv"
  `include "output_controller.sv"
  `include "assertion_reporter.sv"
  `include "signal_reporter.sv"
  `include "monitor.sv"
  `include "transaction_table.sv"
  `include "lfsr.sv"
  `include "lfsr_1.sv"
endpackage : sv_basic_comp_pkg
