--
-- TESTBENCH.vhd: fl_extract testbench
-- Copyright (C) 2007 CESNET
-- Author(s): Vlastimil Kosar <xkosar02@stud.fit.vutbr.cz>
--
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above copyright
--    notice, this list of conditions and the following disclaimer in
--    the documentation and/or other materials provided with the
--    distribution.
-- 3. Neither the name of the Company nor the names of its contributors
--    may be used to endorse or promote products derived from this
--    software without specific prior written permission.
--
-- This software is provided ``as is'', and any express or implied
-- warranties, including, but not limited to, the implied warranties of
-- merchantability and fitness for a particular purpose are disclaimed.
-- In no event shall the company or contributors be liable for any
-- direct, indirect, incidental, special, exemplary, or consequential
-- damages (including, but not limited to, procurement of substitute
-- goods or services; loss of use, data, or profits; or business
-- interruption) however caused and on any theory of liability, whether
-- in contract, strict liability, or tort (including negligence or
-- otherwise) arising in any way out of the use of this software, even
-- if advised of the possibility of such damage.
--
-- $Id$
--
-- TODO:
--
--
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_textio.all;
use ieee.numeric_std.all;
use std.textio.all;
use work.fl_pkg.all; 
use work.fl_sim_oper.all; 

-- ----------------------------------------------------------------------------
--                        Entity declaration
-- ----------------------------------------------------------------------------
entity TESTBENCH is
end entity TESTBENCH;

-- ----------------------------------------------------------------------------
--                      Architecture declaration
-- ----------------------------------------------------------------------------
architecture TESTBENCH_arch of TESTBENCH is


-- -----------------------Testbench constant-----------------------------------
   constant clkper_50       : time := 20 ns;
   constant clkper_100      : time := 10 ns;
   constant reset_time      : time := 100 * clkper_100;
   constant TX_DATA_WIDTH_X : integer   := 32;

   constant DATA_WIDTH : integer := 32;
   constant PIPELINE_EN: boolean := false;
   constant PACKET_NO: integer := 1;
   constant OFFSET: integer := 4;
   constant SIZE: integer := 15;
-- -----------------------Testbench auxilarity signals-------------------------
     -- CLK_GEN Signals
     signal reset             : std_logic;
     signal clk               : std_logic;
     signal clk_50_in         : std_logic;
     signal clk50             : std_logic;
     signal clk100            : std_logic;
     signal lock              : std_logic;
     signal fl_clk            : std_logic;

     -- Frame Link Bus 32 (FL_SIM)
     signal FL_bus    : t_fl32;
     signal OUT_BUS   : t_fl32;
   
     -- FL_SIM component ctrl      
     signal fl_sim_ctrl        : t_fl_ctrl;
     signal fl_sim_strobe      : std_logic;
     signal fl_sim_busy        : std_logic;

     signal EXT_DATA : std_logic_vector(SIZE*8-1 downto 0);
     signal EXT_DATA_VLD : std_logic;
     
begin

-- Reset generation -----------------------------------------------------------
   reset_gen : process
   begin
      reset <= '1';
      wait for reset_time;
      reset <= '0';
      wait;
   end process reset_gen;
   
-- clk50 generator ------------------------------------------------------------
clk50_gen : process
begin
   clk_50_in <= '1';
   wait for clkper_50/2;
   clk_50_in <= '0';
   wait for clkper_50/2;
end process;

-- CLK_GEN component ----------------------------------------------------------
CLK_GEN_U: entity work.CLK_GEN
   port map (
      -- Input
      CLK50_IN    => clk_50_in,
      RESET       => '0',
      -- Output
      CLK50_OUT   => clk50,
      CLK25       => open,
      CLK100      => clk100,
      CLK200      => open,
      LOCK        => lock
   );
clk <= clk100;
fl_clk <= clk100;

-- Frame Link Bus simulation component ------------------------------------------
FL_SIM_U : entity work.FL_SIM
   generic map (
      DATA_WIDTH=>TX_DATA_WIDTH_X,
      FRAME_PARTS => 3
   )
   port map (
      -- Common interface
      FL_RESET           => reset,
      FL_CLK             => fl_clk,

      -- FL Bus Interface
      RX_DATA=>(others => '0'),
      RX_REM=>(others => '0'),
      RX_SOF_N=>'1',
      RX_EOF_N=>'1',
      RX_SOP_N=>'1',
      RX_EOP_N=>'1',
      RX_SRC_RDY_N=>'1',
      RX_DST_RDY_N=>open,

      TX_DATA=>FL_bus.DATA,
      TX_REM=>FL_bus.DREM,
      TX_SOF_N=>FL_bus.SOF_N,
      TX_EOF_N=>FL_bus.EOF_N,
      TX_SOP_N=>FL_bus.SOP_N,
      TX_EOP_N=>FL_bus.EOP_N,
      TX_SRC_RDY_N=>FL_bus.SRC_RDY_N,
      TX_DST_RDY_N=>FL_bus.DST_RDY_N,

      -- IB SIM interface
      CTRL               => fl_sim_ctrl,
      STROBE             => fl_sim_strobe,
      BUSY               => fl_sim_busy
     );

FL_EXTRACT_U: entity work.FL_EXTRACT
  generic map(
      -- Frame link width
      DATA_WIDTH=>DATA_WIDTH,
      PIPELINE_EN=>PIPELINE_EN, -- Enable registers on output fl interface

      -- Header / Footer data present
      PACKET_NO=>PACKET_NO, -- Part of Frame where the field is extracted

      -- Extract option
      OFFSET=>OFFSET, -- Start extracting on specified offset
      SIZE=>SIZE  -- Size of "Extracted field" in Bytes
      )
   port map(
      CLK=>FL_CLK,
      RESET=>RESET,

      EXT_DATA=>EXT_DATA,
      EXT_DATA_VLD=>EXT_DATA_VLD,

      -- Input Interface
      RX_DATA=>FL_bus.DATA,
      RX_REM=>FL_bus.DREM,
      RX_SRC_RDY_N=>FL_bus.SRC_RDY_N,
      RX_DST_RDY_N=>FL_bus.DST_RDY_N,
      RX_SOP_N=>FL_bus.SOP_N,
      RX_EOP_N=>FL_bus.EOP_N,
      RX_SOF_N=>FL_bus.SOF_N,
      RX_EOF_N=>FL_bus.EOF_N,

      -- Output Interface
      TX_DATA=>OUT_BUS.DATA,
      TX_REM=>OUT_BUS.DREM,
      TX_SRC_RDY_N=>OUT_BUS.SRC_RDY_N,
      TX_DST_RDY_N=>OUT_BUS.DST_RDY_N,
      TX_SOP_N=>OUT_BUS.SOP_N,
      TX_EOP_N=>OUT_BUS.EOP_N,
      TX_SOF_N=>OUT_BUS.SOF_N,
      TX_EOF_N=>OUT_BUS.EOF_N
   );

OUT_BUS.DST_RDY_N<='0';

tb : process
-- support function
procedure fl_op(ctrl : in t_fl_ctrl) is
begin
   wait until (FL_CLK'event and FL_CLK='1' and fl_sim_busy = '0');
   fl_sim_ctrl <= ctrl;
   fl_sim_strobe <= '1';
   wait until (FL_CLK'event and FL_CLK='1');
   fl_sim_strobe <= '0';
end fl_op;

begin
-- Testbench
fl_sim_strobe <= '0';
wait for reset_time;
fl_op(fl_send32("../../../debug/sim/sim/tests/fl_sim.txt"));
fl_op(fl_send32("../../../debug/sim/sim/tests/fl_sim2.txt"));
end process;
end architecture TESTBENCH_arch;
