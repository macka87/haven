/* *****************************************************************************
 * Project Name: Genetic Algorithm for ALU
 * File Name:    sv_alu_coverage_pkg.sv
 * Description:  UVM Genetic Algorithm Components Package.
 * Authors:      Marcela Simkova <isimkova@fit.vutbr.cz> 
 * Date:         13.2.2014
 * ************************************************************************** */

 package sv_alu_coverage_pkg; 
  
   // Includes
   `include "alu_coverage_info.svh"
   
 endpackage : sv_alu_coverage_pkg
