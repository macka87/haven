--
-- ib_switch_mux.vhd: ib_switch output multiplexor
-- Copyright (C) 2006 CESNET
-- Author(s): Petr Kobiersky <xkobie00@stud.fit.vutbr.cz>
--            Patrik Beck <beck@liberouter.org>
--
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above copyright
--    notice, this list of conditions and the following disclaimer in
--    the documentation and/or other materials provided with the
--    distribution.
-- 3. Neither the name of the Company nor the names of its contributors
--    may be used to endorse or promote products derived from this
--    software without specific prior written permission.
--
-- This software is provided ``as is'', and any express or implied
-- warranties, including, but not limited to, the implied warranties of
-- merchantability and fitness for a particular purpose are disclaimed.
-- In no event shall the company or contributors be liable for any
-- direct, indirect, incidental, special, exemplary, or consequential
-- damages (including, but not limited to, procurement of substitute
-- goods or services; loss of use, data, or profits; or business
-- interruption) however caused and on any theory of liability, whether
-- in contract, strict liability, or tort (including negligence or
-- otherwise) arising in any way out of the use of this software, even
-- if advised of the possibility of such damage.
--
-- $Id$
--
-- TODO:
--
--
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use work.math_pack.all;
-- ----------------------------------------------------------------------------
--                        Entity declaration
-- ----------------------------------------------------------------------------
entity CB_SWITCH_MUX is
   generic(
      DATA_WIDTH  :  INTEGER := 16;
      DS_PORTS    :  INTEGER := 2
   );
   port(
   
   -- Upstream
   PORT0_DATA_IN  : in std_logic_vector(DATA_WIDTH-1 downto 0);
   PORT0_DATA_OUT : out std_logic_vector(DATA_WIDTH-1 downto 0);

   -- Downstream
   DS_DATA_IN  : in std_logic_vector((DS_PORTS*DATA_WIDTH)-1 downto 0);
   DS_DATA_OUT : out std_logic_vector((DS_PORTS*DATA_WIDTH)-1 downto 0);
  
   PORT0_MUX_SEL  : in std_logic_vector(LOG2(DS_PORTS)-1 downto 0)
  
   );
end entity CB_SWITCH_MUX;

-- ----------------------------------------------------------------------------
--                      Architecture declaration
-- ----------------------------------------------------------------------------
architecture CB_SWITCH_MUX_ARCH of CB_SWITCH_MUX is


begin

-- multiplexor port0 ----------------------------------------------------------
process(PORT0_MUX_SEL, DS_DATA_IN)
begin
   PORT0_DATA_OUT <= DS_DATA_IN(DATA_WIDTH-1 downto 0);
   for i in 0 to DS_PORTS-1 loop
      if(conv_std_logic_vector(i, LOG2(DS_PORTS)) = PORT0_MUX_SEL) then
         PORT0_DATA_OUT <= DS_DATA_IN((DATA_WIDTH*(i + 1))-1 downto DATA_WIDTH*i);
      end if;
   end loop;
end process;
                              
OUT_G: for i in 0 to DS_PORTS-1 generate
   DS_DATA_OUT((i+1)*DATA_WIDTH-1 downto i*DATA_WIDTH) <= PORT0_DATA_IN;
end generate;

end architecture CB_SWITCH_MUX_ARCH;

