--
-- comparator.vhd : </=/> comparator
-- Copyright (C) 2008 CESNET
-- Author(s): Tomas Malek <tomalek@liberouter.org>
--
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above copyright
--    notice, this list of conditions and the following disclaimer in
--    the documentation and/or other materials provided with the
--    distribution.
-- 3. Neither the name of the Company nor the names of its contributors
--    may be used to endorse or promote products derived from this
--    software without specific prior written permission.
--
-- This software is provided ``as is'', and any express or implied
-- warranties, including, but not limited to, the implied warranties of
-- merchantability and fitness for a particular purpose are disclaimed.
-- In no event shall the company or contributors be liable for any
-- direct, indirect, incidental, special, exemplary, or consequential
-- damages (including, but not limited to, procurement of substitute
-- goods or services; loss of use, data, or profits; or business
-- interruption) however caused and on any theory of liability, whether
-- in contract, strict liability, or tort (including negligence or
-- otherwise) arising in any way out of the use of this software, even
-- if advised of the possibility of such damage.
--
-- $Id$
--
-- TODO:
--

library IEEE;  
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;

library unisim;
use unisim.vcomponents.all;

-- ----------------------------------------------------------------------------
--                   ENTITY DECLARATION -- </=/> comparator                  -- 
-- ----------------------------------------------------------------------------

entity COMPARATOR is 
   generic(
      WIDTH   : integer:= 64
   ); 
   port (

      -- Input interface ------------------------------------------------------
      ADDR  : in  std_logic_vector(WIDTH-1 downto 0);
      CONST : in  std_logic_vector(WIDTH-1 downto 0);      

      -- Output interface -----------------------------------------------------
      EQ    : out std_logic;
      LT_GT : out std_logic
   );
end COMPARATOR;

-- ----------------------------------------------------------------------------
--               ARCHITECTURE DECLARATION  --  </=/> comparator              --
-- ----------------------------------------------------------------------------

architecture comparator_arch of COMPARATOR is

   signal sub_result : std_logic_vector(WIDTH downto 0);

begin

   -- -------------------------------------------------------------------------
   --                       SOLUTION USING SUBTRACTER                        --
   -- -------------------------------------------------------------------------

   -- 'ADDR - CONST' substracter ----------------------------------------------
   --sub_resultp: process(ADDR, CONST)
   --begin
   --   sub_result <= ext(ADDR,WIDTH+1) - ext(CONST,WIDTH+1);
   --end process;

   -- 'recognize result' decoder ----------------------------------------------
   --EQ     <=  '1' when sub_result = 0 else 
   --           '0';   
   --            
   --LT_GT  <=  not sub_result(WIDTH);

   -- -------------------------------------------------------------------------
   --                       SOLUTION USING COMPARATORS                       --
   -- -------------------------------------------------------------------------

   process (ADDR, CONST)
   begin
      EQ    <= '0';
      LT_GT <= '0';
      if (ADDR = CONST) then
         EQ <= '1';
      elsif (ADDR > CONST) then
         LT_GT <= '1';
      end if;
   end process;

end comparator_arch;

                     

