/*
 * sv_f2f_pkg.sv: SystemVerilog Fifo2nFifo package
 * Copyright (C) 2008 CESNET
 * Author(s): Marcela Simkova <xsimko03@stud.fit.vutbr.cz>
 *
 * Redistribution and use in source and binary forms, with or without
 * modification, are permitted provided that the following conditions
 * are met:
 * 1. Redistributions of source code must retain the above copyright
 *    notice, this list of conditions and the following disclaimer.
 * 2. Redistributions in binary form must reproduce the above copyright
 *    notice, this list of conditions and the following disclaimer in
 *    the documentation and/or other materials provided with the
 *    distribution.
 * 3. Neither the name of the Company nor the names of its contributors
 *    may be used to endorse or promote products derived from this
 *    software without specific prior written permission.
 *
 * This software is provided ``as is'', and any express or implied
 * warranties, including, but not limited to, the implied warranties of
 * merchantability and fitness for a particular purpose are disclaimed.
 * In no event shall the company or contributors be liable for any
 * direct, indirect, incidental, special, exemplary, or consequential
 * damages (including, but not limited to, procurement of substitute
 * goods or services; loss of use, data, or profits; or business
 * interruption) however caused and on any theory of liability, whether
 * in contract, strict liability, or tort (including negligence or
 * otherwise) arising in any way out of the use of this software, even
 * if advised of the possibility of such damage.
 *
 *
 * TODO:
 */

// Fifo2nFifo Interface
`include "buffer_ifc.sv"

package sv_buffer_pkg; 

  import sv_common_pkg::*; // Import SV common classes

  `include "buffer_transaction.sv"
  `include "fifo_driver.sv"
  `include "nfifo_driver.sv"
  `include "mem_driver.sv"
  `include "fifo_monitor.sv"
  `include "nfifo_monitor.sv"
  `include "mem_monitor.sv"
  `include "mem_monitor_new.sv"
  `include "fifo_responder.sv"
  `include "nfifo_responder.sv"
  `include "mem_responder.sv"
  
endpackage : sv_buffer_pkg
