jbdbgfsy
shfjkghdf