jbdbgfsy