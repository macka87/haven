/* *****************************************************************************
 * Project Name: Genetic Algorithm for ALU
 * File Name:    alu_coverage_info.svh
 * Description:  Information about coverage for ALU.
 * Authors:      Marcela Simkova <isimkova@fit.vutbr.cz> 
 * Date:         13.2.2014
 * ************************************************************************** */

/*!
 * \brief AluCoverageInfo
 * 
 * This class stores information about ALU coverage.
 */
 
 class AluCoverageInfo;
    
  /*! 
   * Data Members
   */  
   
   real alu_in_coverage = 0;
   real alu_out_coverage = 0;
       
 endclass: AluCoverageInfo