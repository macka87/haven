/* *****************************************************************************
 * Project Name: HAVEN - Genetic Algorithm
 * File Name:    sv_alu_coverage_pkg.sv
 * Description:  UVM Genetic Algorithm Components Package.
 * Authors:      Marcela Simkova <isimkova@fit.vutbr.cz> 
 * Date:         2.8.2013
 * ************************************************************************** */

 package sv_alu_coverage_pkg; 
  
   // Standard UVM import & include
   import uvm_pkg::*;
   `include "uvm_macros.svh"
  
   // Includes
   `include "alu_coverage_info.svh"
   
 endpackage : sv_alu_coverage_pkg
