--
-- obuf_gmii_top1_empty.vhd: obuf top level - empty architecture
-- Copyright (C) 2005 CESNET
-- Author(s): Martin Mikusek <martin.mikusek@liberouter.org>
--
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above copyright
--    notice, this list of conditions and the following disclaimer in
--    the documentation and/or other materials provided with the
--    distribution.
-- 3. Neither the name of the Company nor the names of its contributors
--    may be used to endorse or promote products derived from this
--    software without specific prior written permission.
--
-- This software is provided ``as is'', and any express or implied
-- warranties, including, but not limited to, the implied warranties of
-- merchantability and fitness for a particular purpose are disclaimed.
-- In no event shall the company or contributors be liable for any
-- direct, indirect, incidental, special, exemplary, or consequential
-- damages (including, but not limited to, procurement of substitute
-- goods or services; loss of use, data, or profits; or business
-- interruption) however caused and on any theory of liability, whether
-- in contract, strict liability, or tort (including negligence or
-- otherwise) arising in any way out of the use of this software, even
-- if advised of the possibility of such damage.
--
-- $Id$
--
-- TODO:
--
--

----------------------------------------------------------------------------
--                      Architecture declaration
----------------------------------------------------------------------------
architecture empty of obuf_gmii_top1 is

signal empty_sig : std_logic_vector(3 + ((DATA_PATHS*8) + (log2(DATA_PATHS))+5) + 21 - 1 downto 0);
begin
   empty_sig <= RESET   &
                WRCLK   &  -- 3
          		 REFCLK   &

               DATA        &
               DREM        &
               SRC_RDY_N   &
               SOF_N       &
               SOP_N       &
               EOF_N       &
               EOP_N       &

               LBCLK   &
		         LBFRAME &
               LBAS    &  -- 5
               LBRW    &
               LBLAST  &
               LBAD;      --16
      

   TXCLK    <= '0';
   TXD      <= (others => '0');
   TXEN     <= '0';
   TXER     <= '0';
   DST_RDY_N   <= '0';

   LBHOLDA  <= 'Z';
   LBRDY    <= 'Z';
   LBAD     <= (others => 'Z');

end architecture empty;

