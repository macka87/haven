/* *****************************************************************************
 * Project Name: Genetic Algorithm for ALU
 * File Name:    chromosome_array.svh
 * Description:  Array of chromosomes.
 * Authors:      Marcela Simkova <isimkova@fit.vutbr.cz> 
 * Date:         13.2.2014
 * ************************************************************************** */

/*!
 * \brief ChromosomeArray
 * 
 * This class represents an array of chromosomes.
 */
 
 class AluChromosomeArray;
    
  /*! 
   * Data Members
   */  
   AluChromosome  alu_chromosome[];  // ALU Chromosomes
   
 endclass: AluChromosomeArray
