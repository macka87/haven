package sv_codix_ca_dpi_pkg;

	import ovm_pkg::*;
	import sv_codix_ca_param_pkg::*;
	import sv_codix_ca_seq_pkg::*;
        import dpi_wrapper_pkg::*;

	`include "ovm_macros.svh"
	`include "input_wrapper.sv"
	`include "output_wrapper.sv"

endpackage
