-- fsm_valid.vhd: FrameLink cutter: FSM Valid
-- (extract and optionally remove data on defined offset in defined frame part)
-- Copyright (C) 2008 CESNET
-- Author(s): Bronislav Pribyl <xpriby12@stud.fit.vutbr.cz>
--
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above copyright
--    notice, this list of conditions and the following disclaimer in
--    the documentation and/or other materials provided with the
--    distribution.
-- 3. Neither the name of the Company nor the names of its contributors
--    may be used to endorse or promote products derived from this
--    software without specific prior written permission.
--
-- This software is provided ``as is'', and any express or implied
-- warranties, including, but not limited to, the implied warranties of
-- merchantability and fitness for a particular purpose are disclaimed.
-- In no event shall the company or contributors be liable for any
-- direct, indirect, incidental, special, exemplary, or consequential
-- damages (including, but not limited to, procurement of substitute
-- goods or services; loss of use, data, or profits; or business
-- interruption) however caused and on any theory of liability, whether
-- in contract, strict liability, or tort (including negligence or
-- otherwise) arising in any way out of the use of this software, even
-- if advised of the possibility of such damage.
--
-- $Id$
--


library ieee;
use ieee.std_logic_1164.all;
use work.math_pack.all;

-- ----------------------------------------------------------------------------
--                      Architecture declaration
-- ----------------------------------------------------------------------------
architecture full of fsm_valid is

   -- ============================== TYPES =====================================

   type t_fsm_valid    is (sv_invalid, sv_valid, sv_done);


   -- ============================== SIGNALS ===================================
   
   signal valid_c_state : t_fsm_valid;
   signal valid_n_state : t_fsm_valid;
   
   
begin

   -- current state register
   Valid_fsm_current_state: process(CLK, RESET)
   begin
      if (RESET = '1') then -- asynchronous reset
         valid_c_state <= sv_invalid;
      elsif (CLK'event and CLK ='1') then
         if (SYN_RESET = '1') then -- synchronous reset
            valid_c_state <= sv_invalid;
         else
            valid_c_state <= valid_n_state;
         end if;
      end if;
   end process;


   -- next state logic
   Valid_fsm_next_state:
   process(valid_c_state, CUT_EXTRACTED)
   begin
      valid_n_state <= sv_invalid;

      case valid_c_state is

         -- invalid
         when sv_invalid =>
            if (cut_extracted = '1') then
               valid_n_state <= sv_valid;
            else
               valid_n_state <= sv_invalid;
            end if;

         -- valid
         when sv_valid =>
            valid_n_state <= sv_done;

         -- done
         when sv_done =>
            valid_n_state <= sv_done;

         -- undefined
         when others =>

      end case;
   end process;


   -- output logic
   Valid_fsm_output: process(valid_c_state)
   begin
      CUT_VLD <= '0';

      case valid_c_state is

         -- invalid
         when sv_invalid =>
            CUT_VLD <= '0';

         -- valid
         when sv_valid =>
            CUT_VLD <= '1';

         -- done
         when sv_done =>
            CUT_VLD <= '0';

         -- undefined
         when others =>

      end case;
   end process;

end architecture full;
