-- fl2cmd.vhd: Entity of FrameLink to Command protocol conversion tool.
-- Copyright (C) 2006 CESNET
-- Author(s): Martin Louda <sandin@liberouter.org>
--
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above copyright
--    notice, this list of conditions and the following disclaimer in
--    the documentation and/or other materials provided with the
--    distribution.
-- 3. Neither the name of the Company nor the names of its contributors
--    may be used to endorse or promote products derived from this
--    software without specific prior written permission.
--
-- This software is provided ``as is'', and any express or implied
-- warranties, including, but not limited to, the implied warranties of
-- merchantability and fitness for a particular purpose are disclaimed.
-- In no event shall the company or contributors be liable for any
-- direct, indirect, incidental, special, exemplary, or consequential
-- damages (including, but not limited to, procurement of substitute
-- goods or services; loss of use, data, or profits; or business
-- interruption) however caused and on any theory of liability, whether
-- in contract, strict liability, or tort (including negligence or
-- otherwise) arising in any way out of the use of this software, even
-- if advised of the possibility of such damage.
--
-- $Id$
--
-- TODO:
--

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

-- library containing log2 function
use work.math_pack.all;

-- ------------------------------------------------------------------------
--                        Entity declaration
-- ------------------------------------------------------------------------
entity FL2CMD is
   generic(
      -- FL /CMD data bus width
      -- only 8, 16, 32, 64 and 128 supported
      DATA_WIDTH  : integer;
      -- Header data present
      HEADER      : boolean := true;
      -- Footer data present
      FOOTER      : boolean := true
   );
   port(
      CLK            : in  std_logic;
      RESET          : in  std_logic;

      -- FL interface
      FL_DATA        : in  std_logic_vector(DATA_WIDTH-1 downto 0);
      FL_REM         : in  std_logic_vector(log2(DATA_WIDTH/8)-1 downto 0);
      FL_SOF_N       : in  std_logic;
      FL_EOF_N       : in  std_logic;
      FL_SOP_N       : in  std_logic;
      FL_EOP_N       : in  std_logic;
      FL_SRC_RDY_N   : in  std_logic;
      FL_DST_RDY_N   : out std_logic;

      -- CMD interface
      CMD_DATA       : out std_logic_vector(DATA_WIDTH-1 downto 0);
      CMD_COMMAND    : out std_logic_vector((DATA_WIDTH/8)-1 downto 0);
      CMD_SRC_RDY    : out std_logic;
      CMD_DST_RDY    : in  std_logic
   );
end entity FL2CMD;
