/* *****************************************************************************
 * Project Name: Random Search for ALU
 * File Name:    sv_alu_rs_pkg.sv
 * Description:  Random Search Components Package.
 * Authors:      Marcela Simkova <isimkova@fit.vutbr.cz> 
 * Date:         17.6.2014
 * ************************************************************************** */

 package sv_alu_rs_pkg; 
  
   // Package imports
   import sv_alu_seq_pkg::*;     
   import sv_alu_param_pkg::*;
   import sv_alu_env_pkg::*;
   import sv_alu_ga_pkg::*;
   import sv_alu_coverage_pkg::*;
   
   // Includes
   `include "alu_rs_input_transaction.svh"
   `include "transaction_rs_sequencer.svh"
   `include "alu_rs_agent.svh"
    
 endpackage : sv_alu_rs_pkg
