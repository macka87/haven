/*
 * testbench_8_64.sv: Top Entity for IB_TRANSFORMER automatic test
 * Copyright (C) 2008 CESNET
 * Author(s): Tomas Malek <tomalek@liberouter.org>
 *
 * Redistribution and use in source and binary forms, with or without
 * modification, are permitted provided that the following conditions
 * are met:
 * 1. Redistributions of source code must retain the above copyright
 *    notice, this list of conditions and the following disclaimer.
 * 2. Redistributions in binary form must reproduce the above copyright
 *    notice, this list of conditions and the following disclaimer in
 *    the documentation and/or other materials provided with the
 *    distribution.
 * 3. Neither the name of the Company nor the names of its contributors
 *    may be used to endorse or promote products derived from this
 *    software without specific prior written permission.
 *
 * This software is provided ``as is'', and any express or implied
 * warranties, including, but not limited to, the implied warranties of
 * merchantability and fitness for a particular purpose are disclaimed.
 * In no event shall the company or contributors be liable for any
 * direct, indirect, incidental, special, exemplary, or consequential
 * damages (including, but not limited to, procurement of substitute
 * goods or services; loss of use, data, or profits; or business
 * interruption) however caused and on any theory of liability, whether
 * in contract, strict liability, or tort (including negligence or
 * otherwise) arising in any way out of the use of this software, even
 * if advised of the possibility of such damage.
 *
 * $Id: testbench_8_64.sv 1899 2008-03-26 15:52:13Z tomalek $
 *
 * TODO:
 *
 */
 
import test_pkg::*; // Test constants and types

// ----------------------------------------------------------------------------
//                                 TESTBENCH
// ----------------------------------------------------------------------------
module testbench;

  // -- Testbench wires and registers -----------------------------------------
  logic CLK   = 0;
  logic RESET;

  iIB64 UP_IN      (CLK, RESET);
  iIB64 UP_OUT     (CLK, RESET);
  iIB8  DOWN_OUT   (CLK, RESET);
  iIB8  DOWN_IN    (CLK, RESET);  
  
  //-- Clock generation -------------------------------------------------------
  always #(cClkPeriod/2) CLK = ~CLK;

  //-- Unit Under Test --------------------------------------------------------
  IB_TRANSFORMER_8_64_SV UUT (.CLK          (CLK),
                              .RESET        (RESET),
                              .UP_IN        (UP_IN   ),
                              .UP_OUT       (UP_OUT  ),
                              .DOWN_OUT     (DOWN_OUT),
                              .DOWN_IN      (DOWN_IN )
                             );

  //-- Test -------------------------------------------------------------------
  TEST_8_64 TEST_U           (.CLK          (CLK),
                              .RESET        (RESET),
                              .UP_IN        (UP_IN   ),
                              .UP_OUT       (UP_OUT  ),
                              .DOWN_OUT     (DOWN_OUT),
                              .DOWN_IN      (DOWN_IN )                        
                             );
endmodule : testbench



